library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity tabelas is
	port(
		ENDERECOS_AUDIO : in std_logic_vector(8 downto 0);
		nota				 :	in std_logic_vector(3 downto 0);
		clk				 :	in std_logic;
		DADOS_AUDIO		 : out std_logic_vector(15 downto 0);
		LARGURA_ENDERECOS_AUDIO	: out std_logic_vector(8 downto 0);
		reset				 :	out std_logic
	);end tabelas;
	
architecture behavior of tabelas is
	signal aux_nota : integer range 0 to 12;
	signal aux_dados : integer range 0 to 511;
	signal n_pontos : integer range 0 to 511;
begin

	aux_dados <= to_integer(unsigned(ENDERECOS_AUDIO));
	aux_nota <= to_integer(unsigned(nota));
	LARGURA_ENDERECOS_AUDIO <= std_logic_vector(to_unsigned(n_pontos,9));
	 
	process(clk)
		begin
			case aux_nota is
				when 1 =>
					n_pontos <= 366;
					reset <= '0';
					case aux_dados is
					    when  0  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  1  =>    DADOS_AUDIO <=  "0000001000110100";
						 when  2  =>    DADOS_AUDIO <=  "0000010001100111";
						 when  3  =>    DADOS_AUDIO <=  "0000011010011011";
						 when  4  =>    DADOS_AUDIO <=  "0000100011001110";
						 when  5  =>    DADOS_AUDIO <=  "0000101100000000";
						 when  6  =>    DADOS_AUDIO <=  "0000110100110010";
						 when  7  =>    DADOS_AUDIO <=  "0000111101100010";
						 when  8  =>    DADOS_AUDIO <=  "0001000110010010";
						 when  9  =>    DADOS_AUDIO <=  "0001001111000000";
						 when  10  =>    DADOS_AUDIO <=  "0001010111101100";
						 when  11  =>    DADOS_AUDIO <=  "0001100000010111";
						 when  12  =>    DADOS_AUDIO <=  "0001101001000000";
						 when  13  =>    DADOS_AUDIO <=  "0001110001100111";
						 when  14  =>    DADOS_AUDIO <=  "0001111010001100";
						 when  15  =>    DADOS_AUDIO <=  "0010000010101111";
						 when  16  =>    DADOS_AUDIO <=  "0010001011001111";
						 when  17  =>    DADOS_AUDIO <=  "0010010011101100";
						 when  18  =>    DADOS_AUDIO <=  "0010011100000111";
						 when  19  =>    DADOS_AUDIO <=  "0010100100011111";
						 when  20  =>    DADOS_AUDIO <=  "0010101100110011";
						 when  21  =>    DADOS_AUDIO <=  "0010110101000101";
						 when  22  =>    DADOS_AUDIO <=  "0010111101010011";
						 when  23  =>    DADOS_AUDIO <=  "0011000101011101";
						 when  24  =>    DADOS_AUDIO <=  "0011001101100011";
						 when  25  =>    DADOS_AUDIO <=  "0011010101100110";
						 when  26  =>    DADOS_AUDIO <=  "0011011101100101";
						 when  27  =>    DADOS_AUDIO <=  "0011100101011111";
						 when  28  =>    DADOS_AUDIO <=  "0011101101010101";
						 when  29  =>    DADOS_AUDIO <=  "0011110101000111";
						 when  30  =>    DADOS_AUDIO <=  "0011111100110100";
						 when  31  =>    DADOS_AUDIO <=  "0100000100011100";
						 when  32  =>    DADOS_AUDIO <=  "0100001011111111";
						 when  33  =>    DADOS_AUDIO <=  "0100010011011101";
						 when  34  =>    DADOS_AUDIO <=  "0100011010110110";
						 when  35  =>    DADOS_AUDIO <=  "0100100010001001";
						 when  36  =>    DADOS_AUDIO <=  "0100101001010111";
						 when  37  =>    DADOS_AUDIO <=  "0100110000100000";
						 when  38  =>    DADOS_AUDIO <=  "0100110111100010";
						 when  39  =>    DADOS_AUDIO <=  "0100111110011111";
						 when  40  =>    DADOS_AUDIO <=  "0101000101010101";
						 when  41  =>    DADOS_AUDIO <=  "0101001100000110";
						 when  42  =>    DADOS_AUDIO <=  "0101010010110000";
						 when  43  =>    DADOS_AUDIO <=  "0101011001010100";
						 when  44  =>    DADOS_AUDIO <=  "0101011111110001";
						 when  45  =>    DADOS_AUDIO <=  "0101100110000111";
						 when  46  =>    DADOS_AUDIO <=  "0101101100010111";
						 when  47  =>    DADOS_AUDIO <=  "0101110010100000";
						 when  48  =>    DADOS_AUDIO <=  "0101111000100010";
						 when  49  =>    DADOS_AUDIO <=  "0101111110011100";
						 when  50  =>    DADOS_AUDIO <=  "0110000100010000";
						 when  51  =>    DADOS_AUDIO <=  "0110001001111100";
						 when  52  =>    DADOS_AUDIO <=  "0110001111100000";
						 when  53  =>    DADOS_AUDIO <=  "0110010100111101";
						 when  54  =>    DADOS_AUDIO <=  "0110011010010011";
						 when  55  =>    DADOS_AUDIO <=  "0110011111100000";
						 when  56  =>    DADOS_AUDIO <=  "0110100100100110";
						 when  57  =>    DADOS_AUDIO <=  "0110101001100011";
						 when  58  =>    DADOS_AUDIO <=  "0110101110011001";
						 when  59  =>    DADOS_AUDIO <=  "0110110011000110";
						 when  60  =>    DADOS_AUDIO <=  "0110110111101011";
						 when  61  =>    DADOS_AUDIO <=  "0110111100001000";
						 when  62  =>    DADOS_AUDIO <=  "0111000000011101";
						 when  63  =>    DADOS_AUDIO <=  "0111000100101001";
						 when  64  =>    DADOS_AUDIO <=  "0111001000101100";
						 when  65  =>    DADOS_AUDIO <=  "0111001100100111";
						 when  66  =>    DADOS_AUDIO <=  "0111010000011001";
						 when  67  =>    DADOS_AUDIO <=  "0111010100000010";
						 when  68  =>    DADOS_AUDIO <=  "0111010111100010";
						 when  69  =>    DADOS_AUDIO <=  "0111011010111001";
						 when  70  =>    DADOS_AUDIO <=  "0111011110000111";
						 when  71  =>    DADOS_AUDIO <=  "0111100001001101";
						 when  72  =>    DADOS_AUDIO <=  "0111100100001001";
						 when  73  =>    DADOS_AUDIO <=  "0111100110111100";
						 when  74  =>    DADOS_AUDIO <=  "0111101001100101";
						 when  75  =>    DADOS_AUDIO <=  "0111101100000110";
						 when  76  =>    DADOS_AUDIO <=  "0111101110011101";
						 when  77  =>    DADOS_AUDIO <=  "0111110000101011";
						 when  78  =>    DADOS_AUDIO <=  "0111110010101111";
						 when  79  =>    DADOS_AUDIO <=  "0111110100101010";
						 when  80  =>    DADOS_AUDIO <=  "0111110110011011";
						 when  81  =>    DADOS_AUDIO <=  "0111111000000011";
						 when  82  =>    DADOS_AUDIO <=  "0111111001100001";
						 when  83  =>    DADOS_AUDIO <=  "0111111010110110";
						 when  84  =>    DADOS_AUDIO <=  "0111111100000001";
						 when  85  =>    DADOS_AUDIO <=  "0111111101000010";
						 when  86  =>    DADOS_AUDIO <=  "0111111101111010";
						 when  87  =>    DADOS_AUDIO <=  "0111111110101000";
						 when  88  =>    DADOS_AUDIO <=  "0111111111001100";
						 when  89  =>    DADOS_AUDIO <=  "0111111111100111";
						 when  90  =>    DADOS_AUDIO <=  "0111111111111000";
						 when  91  =>    DADOS_AUDIO <=  "0111111111111111";
						 when  92  =>    DADOS_AUDIO <=  "0111111111111101";
						 when  93  =>    DADOS_AUDIO <=  "0111111111110001";
						 when  94  =>    DADOS_AUDIO <=  "0111111111011011";
						 when  95  =>    DADOS_AUDIO <=  "0111111110111011";
						 when  96  =>    DADOS_AUDIO <=  "0111111110010010";
						 when  97  =>    DADOS_AUDIO <=  "0111111101011111";
						 when  98  =>    DADOS_AUDIO <=  "0111111100100011";
						 when  99  =>    DADOS_AUDIO <=  "0111111011011100";
						 when  100  =>    DADOS_AUDIO <=  "0111111010001100";
						 when  101  =>    DADOS_AUDIO <=  "0111111000110011";
						 when  102  =>    DADOS_AUDIO <=  "0111110111010000";
						 when  103  =>    DADOS_AUDIO <=  "0111110101100011";
						 when  104  =>    DADOS_AUDIO <=  "0111110011101101";
						 when  105  =>    DADOS_AUDIO <=  "0111110001101110";
						 when  106  =>    DADOS_AUDIO <=  "0111101111100101";
						 when  107  =>    DADOS_AUDIO <=  "0111101101010011";
						 when  108  =>    DADOS_AUDIO <=  "0111101010110111";
						 when  109  =>    DADOS_AUDIO <=  "0111101000010010";
						 when  110  =>    DADOS_AUDIO <=  "0111100101100011";
						 when  111  =>    DADOS_AUDIO <=  "0111100010101100";
						 when  112  =>    DADOS_AUDIO <=  "0111011111101011";
						 when  113  =>    DADOS_AUDIO <=  "0111011100100001";
						 when  114  =>    DADOS_AUDIO <=  "0111011001001111";
						 when  115  =>    DADOS_AUDIO <=  "0111010101110011";
						 when  116  =>    DADOS_AUDIO <=  "0111010010001110";
						 when  117  =>    DADOS_AUDIO <=  "0111001110100001";
						 when  118  =>    DADOS_AUDIO <=  "0111001010101010";
						 when  119  =>    DADOS_AUDIO <=  "0111000110101011";
						 when  120  =>    DADOS_AUDIO <=  "0111000010100100";
						 when  121  =>    DADOS_AUDIO <=  "0110111110010100";
						 when  122  =>    DADOS_AUDIO <=  "0110111001111011";
						 when  123  =>    DADOS_AUDIO <=  "0110110101011010";
						 when  124  =>    DADOS_AUDIO <=  "0110110000110001";
						 when  125  =>    DADOS_AUDIO <=  "0110101011111111";
						 when  126  =>    DADOS_AUDIO <=  "0110100111000101";
						 when  127  =>    DADOS_AUDIO <=  "0110100010000100";
						 when  128  =>    DADOS_AUDIO <=  "0110011100111010";
						 when  129  =>    DADOS_AUDIO <=  "0110010111101001";
						 when  130  =>    DADOS_AUDIO <=  "0110010010010000";
						 when  131  =>    DADOS_AUDIO <=  "0110001100101111";
						 when  132  =>    DADOS_AUDIO <=  "0110000111000111";
						 when  133  =>    DADOS_AUDIO <=  "0110000001010111";
						 when  134  =>    DADOS_AUDIO <=  "0101111011100000";
						 when  135  =>    DADOS_AUDIO <=  "0101110101100010";
						 when  136  =>    DADOS_AUDIO <=  "0101101111011100";
						 when  137  =>    DADOS_AUDIO <=  "0101101001010000";
						 when  138  =>    DADOS_AUDIO <=  "0101100010111101";
						 when  139  =>    DADOS_AUDIO <=  "0101011100100011";
						 when  140  =>    DADOS_AUDIO <=  "0101010110000011";
						 when  141  =>    DADOS_AUDIO <=  "0101001111011100";
						 when  142  =>    DADOS_AUDIO <=  "0101001000101110";
						 when  143  =>    DADOS_AUDIO <=  "0101000001111011";
						 when  144  =>    DADOS_AUDIO <=  "0100111011000001";
						 when  145  =>    DADOS_AUDIO <=  "0100110100000010";
						 when  146  =>    DADOS_AUDIO <=  "0100101100111100";
						 when  147  =>    DADOS_AUDIO <=  "0100100101110001";
						 when  148  =>    DADOS_AUDIO <=  "0100011110100000";
						 when  149  =>    DADOS_AUDIO <=  "0100010111001010";
						 when  150  =>    DADOS_AUDIO <=  "0100001111101110";
						 when  151  =>    DADOS_AUDIO <=  "0100001000001110";
						 when  152  =>    DADOS_AUDIO <=  "0100000000101000";
						 when  153  =>    DADOS_AUDIO <=  "0011111000111110";
						 when  154  =>    DADOS_AUDIO <=  "0011110001001110";
						 when  155  =>    DADOS_AUDIO <=  "0011101001011011";
						 when  156  =>    DADOS_AUDIO <=  "0011100001100010";
						 when  157  =>    DADOS_AUDIO <=  "0011011001100110";
						 when  158  =>    DADOS_AUDIO <=  "0011010001100101";
						 when  159  =>    DADOS_AUDIO <=  "0011001001100001";
						 when  160  =>    DADOS_AUDIO <=  "0011000001011000";
						 when  161  =>    DADOS_AUDIO <=  "0010111001001100";
						 when  162  =>    DADOS_AUDIO <=  "0010110000111101";
						 when  163  =>    DADOS_AUDIO <=  "0010101000101010";
						 when  164  =>    DADOS_AUDIO <=  "0010100000010011";
						 when  165  =>    DADOS_AUDIO <=  "0010010111111010";
						 when  166  =>    DADOS_AUDIO <=  "0010001111011110";
						 when  167  =>    DADOS_AUDIO <=  "0010000110111111";
						 when  168  =>    DADOS_AUDIO <=  "0001111110011110";
						 when  169  =>    DADOS_AUDIO <=  "0001110101111010";
						 when  170  =>    DADOS_AUDIO <=  "0001101101010100";
						 when  171  =>    DADOS_AUDIO <=  "0001100100101100";
						 when  172  =>    DADOS_AUDIO <=  "0001011100000010";
						 when  173  =>    DADOS_AUDIO <=  "0001010011010110";
						 when  174  =>    DADOS_AUDIO <=  "0001001010101001";
						 when  175  =>    DADOS_AUDIO <=  "0001000001111010";
						 when  176  =>    DADOS_AUDIO <=  "0000111001001010";
						 when  177  =>    DADOS_AUDIO <=  "0000110000011001";
						 when  178  =>    DADOS_AUDIO <=  "0000100111100111";
						 when  179  =>    DADOS_AUDIO <=  "0000011110110101";
						 when  180  =>    DADOS_AUDIO <=  "0000010110000001";
						 when  181  =>    DADOS_AUDIO <=  "0000001101001110";
						 when  182  =>    DADOS_AUDIO <=  "0000000100011010";
						 when  183  =>    DADOS_AUDIO <=  "1111111011100110";
						 when  184  =>    DADOS_AUDIO <=  "1111110010110010";
						 when  185  =>    DADOS_AUDIO <=  "1111101001111111";
						 when  186  =>    DADOS_AUDIO <=  "1111100001001011";
						 when  187  =>    DADOS_AUDIO <=  "1111011000011001";
						 when  188  =>    DADOS_AUDIO <=  "1111001111100111";
						 when  189  =>    DADOS_AUDIO <=  "1111000110110110";
						 when  190  =>    DADOS_AUDIO <=  "1110111110000110";
						 when  191  =>    DADOS_AUDIO <=  "1110110101010111";
						 when  192  =>    DADOS_AUDIO <=  "1110101100101010";
						 when  193  =>    DADOS_AUDIO <=  "1110100011111110";
						 when  194  =>    DADOS_AUDIO <=  "1110011011010100";
						 when  195  =>    DADOS_AUDIO <=  "1110010010101100";
						 when  196  =>    DADOS_AUDIO <=  "1110001010000110";
						 when  197  =>    DADOS_AUDIO <=  "1110000001100010";
						 when  198  =>    DADOS_AUDIO <=  "1101111001000001";
						 when  199  =>    DADOS_AUDIO <=  "1101110000100010";
						 when  200  =>    DADOS_AUDIO <=  "1101101000000110";
						 when  201  =>    DADOS_AUDIO <=  "1101011111101101";
						 when  202  =>    DADOS_AUDIO <=  "1101010111010110";
						 when  203  =>    DADOS_AUDIO <=  "1101001111000011";
						 when  204  =>    DADOS_AUDIO <=  "1101000110110100";
						 when  205  =>    DADOS_AUDIO <=  "1100111110101000";
						 when  206  =>    DADOS_AUDIO <=  "1100110110011111";
						 when  207  =>    DADOS_AUDIO <=  "1100101110011011";
						 when  208  =>    DADOS_AUDIO <=  "1100100110011010";
						 when  209  =>    DADOS_AUDIO <=  "1100011110011110";
						 when  210  =>    DADOS_AUDIO <=  "1100010110100101";
						 when  211  =>    DADOS_AUDIO <=  "1100001110110010";
						 when  212  =>    DADOS_AUDIO <=  "1100000111000010";
						 when  213  =>    DADOS_AUDIO <=  "1011111111011000";
						 when  214  =>    DADOS_AUDIO <=  "1011110111110010";
						 when  215  =>    DADOS_AUDIO <=  "1011110000010010";
						 when  216  =>    DADOS_AUDIO <=  "1011101000110110";
						 when  217  =>    DADOS_AUDIO <=  "1011100001100000";
						 when  218  =>    DADOS_AUDIO <=  "1011011010001111";
						 when  219  =>    DADOS_AUDIO <=  "1011010011000100";
						 when  220  =>    DADOS_AUDIO <=  "1011001011111110";
						 when  221  =>    DADOS_AUDIO <=  "1011000100111111";
						 when  222  =>    DADOS_AUDIO <=  "1010111110000101";
						 when  223  =>    DADOS_AUDIO <=  "1010110111010010";
						 when  224  =>    DADOS_AUDIO <=  "1010110000100100";
						 when  225  =>    DADOS_AUDIO <=  "1010101001111101";
						 when  226  =>    DADOS_AUDIO <=  "1010100011011101";
						 when  227  =>    DADOS_AUDIO <=  "1010011101000011";
						 when  228  =>    DADOS_AUDIO <=  "1010010110110000";
						 when  229  =>    DADOS_AUDIO <=  "1010010000100100";
						 when  230  =>    DADOS_AUDIO <=  "1010001010011110";
						 when  231  =>    DADOS_AUDIO <=  "1010000100100000";
						 when  232  =>    DADOS_AUDIO <=  "1001111110101001";
						 when  233  =>    DADOS_AUDIO <=  "1001111000111001";
						 when  234  =>    DADOS_AUDIO <=  "1001110011010001";
						 when  235  =>    DADOS_AUDIO <=  "1001101101110000";
						 when  236  =>    DADOS_AUDIO <=  "1001101000010111";
						 when  237  =>    DADOS_AUDIO <=  "1001100011000110";
						 when  238  =>    DADOS_AUDIO <=  "1001011101111100";
						 when  239  =>    DADOS_AUDIO <=  "1001011000111011";
						 when  240  =>    DADOS_AUDIO <=  "1001010100000001";
						 when  241  =>    DADOS_AUDIO <=  "1001001111001111";
						 when  242  =>    DADOS_AUDIO <=  "1001001010100110";
						 when  243  =>    DADOS_AUDIO <=  "1001000110000101";
						 when  244  =>    DADOS_AUDIO <=  "1001000001101100";
						 when  245  =>    DADOS_AUDIO <=  "1000111101011100";
						 when  246  =>    DADOS_AUDIO <=  "1000111001010101";
						 when  247  =>    DADOS_AUDIO <=  "1000110101010110";
						 when  248  =>    DADOS_AUDIO <=  "1000110001011111";
						 when  249  =>    DADOS_AUDIO <=  "1000101101110010";
						 when  250  =>    DADOS_AUDIO <=  "1000101010001101";
						 when  251  =>    DADOS_AUDIO <=  "1000100110110001";
						 when  252  =>    DADOS_AUDIO <=  "1000100011011111";
						 when  253  =>    DADOS_AUDIO <=  "1000100000010101";
						 when  254  =>    DADOS_AUDIO <=  "1000011101010100";
						 when  255  =>    DADOS_AUDIO <=  "1000011010011101";
						 when  256  =>    DADOS_AUDIO <=  "1000010111101110";
						 when  257  =>    DADOS_AUDIO <=  "1000010101001001";
						 when  258  =>    DADOS_AUDIO <=  "1000010010101101";
						 when  259  =>    DADOS_AUDIO <=  "1000010000011011";
						 when  260  =>    DADOS_AUDIO <=  "1000001110010010";
						 when  261  =>    DADOS_AUDIO <=  "1000001100010011";
						 when  262  =>    DADOS_AUDIO <=  "1000001010011101";
						 when  263  =>    DADOS_AUDIO <=  "1000001000110000";
						 when  264  =>    DADOS_AUDIO <=  "1000000111001101";
						 when  265  =>    DADOS_AUDIO <=  "1000000101110100";
						 when  266  =>    DADOS_AUDIO <=  "1000000100100100";
						 when  267  =>    DADOS_AUDIO <=  "1000000011011101";
						 when  268  =>    DADOS_AUDIO <=  "1000000010100001";
						 when  269  =>    DADOS_AUDIO <=  "1000000001101110";
						 when  270  =>    DADOS_AUDIO <=  "1000000001000101";
						 when  271  =>    DADOS_AUDIO <=  "1000000000100101";
						 when  272  =>    DADOS_AUDIO <=  "1000000000001111";
						 when  273  =>    DADOS_AUDIO <=  "1000000000000011";
						 when  274  =>    DADOS_AUDIO <=  "1000000000000001";
						 when  275  =>    DADOS_AUDIO <=  "1000000000001000";
						 when  276  =>    DADOS_AUDIO <=  "1000000000011001";
						 when  277  =>    DADOS_AUDIO <=  "1000000000110100";
						 when  278  =>    DADOS_AUDIO <=  "1000000001011000";
						 when  279  =>    DADOS_AUDIO <=  "1000000010000110";
						 when  280  =>    DADOS_AUDIO <=  "1000000010111110";
						 when  281  =>    DADOS_AUDIO <=  "1000000011111111";
						 when  282  =>    DADOS_AUDIO <=  "1000000101001010";
						 when  283  =>    DADOS_AUDIO <=  "1000000110011111";
						 when  284  =>    DADOS_AUDIO <=  "1000000111111101";
						 when  285  =>    DADOS_AUDIO <=  "1000001001100101";
						 when  286  =>    DADOS_AUDIO <=  "1000001011010110";
						 when  287  =>    DADOS_AUDIO <=  "1000001101010001";
						 when  288  =>    DADOS_AUDIO <=  "1000001111010101";
						 when  289  =>    DADOS_AUDIO <=  "1000010001100011";
						 when  290  =>    DADOS_AUDIO <=  "1000010011111010";
						 when  291  =>    DADOS_AUDIO <=  "1000010110011011";
						 when  292  =>    DADOS_AUDIO <=  "1000011001000100";
						 when  293  =>    DADOS_AUDIO <=  "1000011011110111";
						 when  294  =>    DADOS_AUDIO <=  "1000011110110011";
						 when  295  =>    DADOS_AUDIO <=  "1000100001111001";
						 when  296  =>    DADOS_AUDIO <=  "1000100101000111";
						 when  297  =>    DADOS_AUDIO <=  "1000101000011110";
						 when  298  =>    DADOS_AUDIO <=  "1000101011111110";
						 when  299  =>    DADOS_AUDIO <=  "1000101111100111";
						 when  300  =>    DADOS_AUDIO <=  "1000110011011001";
						 when  301  =>    DADOS_AUDIO <=  "1000110111010100";
						 when  302  =>    DADOS_AUDIO <=  "1000111011010111";
						 when  303  =>    DADOS_AUDIO <=  "1000111111100011";
						 when  304  =>    DADOS_AUDIO <=  "1001000011111000";
						 when  305  =>    DADOS_AUDIO <=  "1001001000010101";
						 when  306  =>    DADOS_AUDIO <=  "1001001100111010";
						 when  307  =>    DADOS_AUDIO <=  "1001010001100111";
						 when  308  =>    DADOS_AUDIO <=  "1001010110011101";
						 when  309  =>    DADOS_AUDIO <=  "1001011011011010";
						 when  310  =>    DADOS_AUDIO <=  "1001100000100000";
						 when  311  =>    DADOS_AUDIO <=  "1001100101101101";
						 when  312  =>    DADOS_AUDIO <=  "1001101011000011";
						 when  313  =>    DADOS_AUDIO <=  "1001110000100000";
						 when  314  =>    DADOS_AUDIO <=  "1001110110000100";
						 when  315  =>    DADOS_AUDIO <=  "1001111011110000";
						 when  316  =>    DADOS_AUDIO <=  "1010000001100100";
						 when  317  =>    DADOS_AUDIO <=  "1010000111011110";
						 when  318  =>    DADOS_AUDIO <=  "1010001101100000";
						 when  319  =>    DADOS_AUDIO <=  "1010010011101001";
						 when  320  =>    DADOS_AUDIO <=  "1010011001111001";
						 when  321  =>    DADOS_AUDIO <=  "1010100000001111";
						 when  322  =>    DADOS_AUDIO <=  "1010100110101100";
						 when  323  =>    DADOS_AUDIO <=  "1010101101010000";
						 when  324  =>    DADOS_AUDIO <=  "1010110011111010";
						 when  325  =>    DADOS_AUDIO <=  "1010111010101011";
						 when  326  =>    DADOS_AUDIO <=  "1011000001100001";
						 when  327  =>    DADOS_AUDIO <=  "1011001000011110";
						 when  328  =>    DADOS_AUDIO <=  "1011001111100000";
						 when  329  =>    DADOS_AUDIO <=  "1011010110101001";
						 when  330  =>    DADOS_AUDIO <=  "1011011101110111";
						 when  331  =>    DADOS_AUDIO <=  "1011100101001010";
						 when  332  =>    DADOS_AUDIO <=  "1011101100100011";
						 when  333  =>    DADOS_AUDIO <=  "1011110100000001";
						 when  334  =>    DADOS_AUDIO <=  "1011111011100100";
						 when  335  =>    DADOS_AUDIO <=  "1100000011001100";
						 when  336  =>    DADOS_AUDIO <=  "1100001010111001";
						 when  337  =>    DADOS_AUDIO <=  "1100010010101011";
						 when  338  =>    DADOS_AUDIO <=  "1100011010100001";
						 when  339  =>    DADOS_AUDIO <=  "1100100010011011";
						 when  340  =>    DADOS_AUDIO <=  "1100101010011010";
						 when  341  =>    DADOS_AUDIO <=  "1100110010011101";
						 when  342  =>    DADOS_AUDIO <=  "1100111010100011";
						 when  343  =>    DADOS_AUDIO <=  "1101000010101101";
						 when  344  =>    DADOS_AUDIO <=  "1101001010111011";
						 when  345  =>    DADOS_AUDIO <=  "1101010011001101";
						 when  346  =>    DADOS_AUDIO <=  "1101011011100001";
						 when  347  =>    DADOS_AUDIO <=  "1101100011111001";
						 when  348  =>    DADOS_AUDIO <=  "1101101100010100";
						 when  349  =>    DADOS_AUDIO <=  "1101110100110001";
						 when  350  =>    DADOS_AUDIO <=  "1101111101010001";
						 when  351  =>    DADOS_AUDIO <=  "1110000101110100";
						 when  352  =>    DADOS_AUDIO <=  "1110001110011001";
						 when  353  =>    DADOS_AUDIO <=  "1110010111000000";
						 when  354  =>    DADOS_AUDIO <=  "1110011111101001";
						 when  355  =>    DADOS_AUDIO <=  "1110101000010100";
						 when  356  =>    DADOS_AUDIO <=  "1110110001000000";
						 when  357  =>    DADOS_AUDIO <=  "1110111001101110";
						 when  358  =>    DADOS_AUDIO <=  "1111000010011110";
						 when  359  =>    DADOS_AUDIO <=  "1111001011001110";
						 when  360  =>    DADOS_AUDIO <=  "1111010100000000";
						 when  361  =>    DADOS_AUDIO <=  "1111011100110010";
						 when  362  =>    DADOS_AUDIO <=  "1111100101100101";
						 when  363  =>    DADOS_AUDIO <=  "1111101110011001";
						 when  364  =>    DADOS_AUDIO <=  "1111110111001100";
						 when  365  =>    DADOS_AUDIO <=  "0000000000000000";
						 when others =>	DADOS_AUDIO <=  "0000000000000000";
					end case;
				when 2 =>
					n_pontos <= 346;
					reset <= '0';
					case aux_dados is
					    when  0  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  1  =>    DADOS_AUDIO <=  "0000001001010100";
						 when  2  =>    DADOS_AUDIO <=  "0000010010101001";
						 when  3  =>    DADOS_AUDIO <=  "0000011011111101";
						 when  4  =>    DADOS_AUDIO <=  "0000100101010000";
						 when  5  =>    DADOS_AUDIO <=  "0000101110100011";
						 when  6  =>    DADOS_AUDIO <=  "0000110111110101";
						 when  7  =>    DADOS_AUDIO <=  "0001000001000110";
						 when  8  =>    DADOS_AUDIO <=  "0001001010010101";
						 when  9  =>    DADOS_AUDIO <=  "0001010011100010";
						 when  10  =>    DADOS_AUDIO <=  "0001011100101110";
						 when  11  =>    DADOS_AUDIO <=  "0001100101111000";
						 when  12  =>    DADOS_AUDIO <=  "0001101111000000";
						 when  13  =>    DADOS_AUDIO <=  "0001111000000101";
						 when  14  =>    DADOS_AUDIO <=  "0010000001001000";
						 when  15  =>    DADOS_AUDIO <=  "0010001010001000";
						 when  16  =>    DADOS_AUDIO <=  "0010010011000101";
						 when  17  =>    DADOS_AUDIO <=  "0010011011111111";
						 when  18  =>    DADOS_AUDIO <=  "0010100100110110";
						 when  19  =>    DADOS_AUDIO <=  "0010101101101001";
						 when  20  =>    DADOS_AUDIO <=  "0010110110011001";
						 when  21  =>    DADOS_AUDIO <=  "0010111111000100";
						 when  22  =>    DADOS_AUDIO <=  "0011000111101100";
						 when  23  =>    DADOS_AUDIO <=  "0011010000001111";
						 when  24  =>    DADOS_AUDIO <=  "0011011000101110";
						 when  25  =>    DADOS_AUDIO <=  "0011100001001001";
						 when  26  =>    DADOS_AUDIO <=  "0011101001011110";
						 when  27  =>    DADOS_AUDIO <=  "0011110001101111";
						 when  28  =>    DADOS_AUDIO <=  "0011111001111010";
						 when  29  =>    DADOS_AUDIO <=  "0100000010000001";
						 when  30  =>    DADOS_AUDIO <=  "0100001010000001";
						 when  31  =>    DADOS_AUDIO <=  "0100010001111100";
						 when  32  =>    DADOS_AUDIO <=  "0100011001110010";
						 when  33  =>    DADOS_AUDIO <=  "0100100001100001";
						 when  34  =>    DADOS_AUDIO <=  "0100101001001010";
						 when  35  =>    DADOS_AUDIO <=  "0100110000101101";
						 when  36  =>    DADOS_AUDIO <=  "0100111000001001";
						 when  37  =>    DADOS_AUDIO <=  "0100111111011111";
						 when  38  =>    DADOS_AUDIO <=  "0101000110101110";
						 when  39  =>    DADOS_AUDIO <=  "0101001101110110";
						 when  40  =>    DADOS_AUDIO <=  "0101010100110110";
						 when  41  =>    DADOS_AUDIO <=  "0101011011110000";
						 when  42  =>    DADOS_AUDIO <=  "0101100010100010";
						 when  43  =>    DADOS_AUDIO <=  "0101101001001101";
						 when  44  =>    DADOS_AUDIO <=  "0101101111110000";
						 when  45  =>    DADOS_AUDIO <=  "0101110110001100";
						 when  46  =>    DADOS_AUDIO <=  "0101111100011111";
						 when  47  =>    DADOS_AUDIO <=  "0110000010101010";
						 when  48  =>    DADOS_AUDIO <=  "0110001000101101";
						 when  49  =>    DADOS_AUDIO <=  "0110001110101000";
						 when  50  =>    DADOS_AUDIO <=  "0110010100011010";
						 when  51  =>    DADOS_AUDIO <=  "0110011010000100";
						 when  52  =>    DADOS_AUDIO <=  "0110011111100101";
						 when  53  =>    DADOS_AUDIO <=  "0110100100111101";
						 when  54  =>    DADOS_AUDIO <=  "0110101010001100";
						 when  55  =>    DADOS_AUDIO <=  "0110101111010010";
						 when  56  =>    DADOS_AUDIO <=  "0110110100001111";
						 when  57  =>    DADOS_AUDIO <=  "0110111001000011";
						 when  58  =>    DADOS_AUDIO <=  "0110111101101101";
						 when  59  =>    DADOS_AUDIO <=  "0111000010001110";
						 when  60  =>    DADOS_AUDIO <=  "0111000110100110";
						 when  61  =>    DADOS_AUDIO <=  "0111001010110011";
						 when  62  =>    DADOS_AUDIO <=  "0111001110110111";
						 when  63  =>    DADOS_AUDIO <=  "0111010010110010";
						 when  64  =>    DADOS_AUDIO <=  "0111010110100010";
						 when  65  =>    DADOS_AUDIO <=  "0111011010001000";
						 when  66  =>    DADOS_AUDIO <=  "0111011101100100";
						 when  67  =>    DADOS_AUDIO <=  "0111100000110110";
						 when  68  =>    DADOS_AUDIO <=  "0111100011111110";
						 when  69  =>    DADOS_AUDIO <=  "0111100110111100";
						 when  70  =>    DADOS_AUDIO <=  "0111101001101111";
						 when  71  =>    DADOS_AUDIO <=  "0111101100011000";
						 when  72  =>    DADOS_AUDIO <=  "0111101110110110";
						 when  73  =>    DADOS_AUDIO <=  "0111110001001010";
						 when  74  =>    DADOS_AUDIO <=  "0111110011010011";
						 when  75  =>    DADOS_AUDIO <=  "0111110101010010";
						 when  76  =>    DADOS_AUDIO <=  "0111110111000110";
						 when  77  =>    DADOS_AUDIO <=  "0111111000110000";
						 when  78  =>    DADOS_AUDIO <=  "0111111010001110";
						 when  79  =>    DADOS_AUDIO <=  "0111111011100010";
						 when  80  =>    DADOS_AUDIO <=  "0111111100101011";
						 when  81  =>    DADOS_AUDIO <=  "0111111101101010";
						 when  82  =>    DADOS_AUDIO <=  "0111111110011101";
						 when  83  =>    DADOS_AUDIO <=  "0111111111000110";
						 when  84  =>    DADOS_AUDIO <=  "0111111111100100";
						 when  85  =>    DADOS_AUDIO <=  "0111111111110111";
						 when  86  =>    DADOS_AUDIO <=  "0111111111111111";
						 when  87  =>    DADOS_AUDIO <=  "0111111111111100";
						 when  88  =>    DADOS_AUDIO <=  "0111111111101111";
						 when  89  =>    DADOS_AUDIO <=  "0111111111010110";
						 when  90  =>    DADOS_AUDIO <=  "0111111110110011";
						 when  91  =>    DADOS_AUDIO <=  "0111111110000101";
						 when  92  =>    DADOS_AUDIO <=  "0111111101001100";
						 when  93  =>    DADOS_AUDIO <=  "0111111100001000";
						 when  94  =>    DADOS_AUDIO <=  "0111111010111010";
						 when  95  =>    DADOS_AUDIO <=  "0111111001100000";
						 when  96  =>    DADOS_AUDIO <=  "0111110111111100";
						 when  97  =>    DADOS_AUDIO <=  "0111110110001110";
						 when  98  =>    DADOS_AUDIO <=  "0111110100010100";
						 when  99  =>    DADOS_AUDIO <=  "0111110010010000";
						 when  100  =>    DADOS_AUDIO <=  "0111110000000001";
						 when  101  =>    DADOS_AUDIO <=  "0111101101101000";
						 when  102  =>    DADOS_AUDIO <=  "0111101011000101";
						 when  103  =>    DADOS_AUDIO <=  "0111101000010111";
						 when  104  =>    DADOS_AUDIO <=  "0111100101011110";
						 when  105  =>    DADOS_AUDIO <=  "0111100010011100";
						 when  106  =>    DADOS_AUDIO <=  "0111011111001111";
						 when  107  =>    DADOS_AUDIO <=  "0111011011110111";
						 when  108  =>    DADOS_AUDIO <=  "0111011000010110";
						 when  109  =>    DADOS_AUDIO <=  "0111010100101011";
						 when  110  =>    DADOS_AUDIO <=  "0111010000110110";
						 when  111  =>    DADOS_AUDIO <=  "0111001100110111";
						 when  112  =>    DADOS_AUDIO <=  "0111001000101110";
						 when  113  =>    DADOS_AUDIO <=  "0111000100011011";
						 when  114  =>    DADOS_AUDIO <=  "0110111111111111";
						 when  115  =>    DADOS_AUDIO <=  "0110111011011001";
						 when  116  =>    DADOS_AUDIO <=  "0110110110101010";
						 when  117  =>    DADOS_AUDIO <=  "0110110001110010";
						 when  118  =>    DADOS_AUDIO <=  "0110101100110000";
						 when  119  =>    DADOS_AUDIO <=  "0110100111100110";
						 when  120  =>    DADOS_AUDIO <=  "0110100010010010";
						 when  121  =>    DADOS_AUDIO <=  "0110011100110101";
						 when  122  =>    DADOS_AUDIO <=  "0110010111010000";
						 when  123  =>    DADOS_AUDIO <=  "0110010001100010";
						 when  124  =>    DADOS_AUDIO <=  "0110001011101100";
						 when  125  =>    DADOS_AUDIO <=  "0110000101101101";
						 when  126  =>    DADOS_AUDIO <=  "0101111111100110";
						 when  127  =>    DADOS_AUDIO <=  "0101111001010110";
						 when  128  =>    DADOS_AUDIO <=  "0101110010111111";
						 when  129  =>    DADOS_AUDIO <=  "0101101100100000";
						 when  130  =>    DADOS_AUDIO <=  "0101100101111001";
						 when  131  =>    DADOS_AUDIO <=  "0101011111001010";
						 when  132  =>    DADOS_AUDIO <=  "0101011000010100";
						 when  133  =>    DADOS_AUDIO <=  "0101010001010111";
						 when  134  =>    DADOS_AUDIO <=  "0101001010010010";
						 when  135  =>    DADOS_AUDIO <=  "0101000011000111";
						 when  136  =>    DADOS_AUDIO <=  "0100111011110101";
						 when  137  =>    DADOS_AUDIO <=  "0100110100011100";
						 when  138  =>    DADOS_AUDIO <=  "0100101100111100";
						 when  139  =>    DADOS_AUDIO <=  "0100100101010110";
						 when  140  =>    DADOS_AUDIO <=  "0100011101101010";
						 when  141  =>    DADOS_AUDIO <=  "0100010101111000";
						 when  142  =>    DADOS_AUDIO <=  "0100001101111111";
						 when  143  =>    DADOS_AUDIO <=  "0100000110000010";
						 when  144  =>    DADOS_AUDIO <=  "0011111101111110";
						 when  145  =>    DADOS_AUDIO <=  "0011110101110101";
						 when  146  =>    DADOS_AUDIO <=  "0011101101100111";
						 when  147  =>    DADOS_AUDIO <=  "0011100101010100";
						 when  148  =>    DADOS_AUDIO <=  "0011011100111100";
						 when  149  =>    DADOS_AUDIO <=  "0011010100011111";
						 when  150  =>    DADOS_AUDIO <=  "0011001011111110";
						 when  151  =>    DADOS_AUDIO <=  "0011000011011001";
						 when  152  =>    DADOS_AUDIO <=  "0010111010101111";
						 when  153  =>    DADOS_AUDIO <=  "0010110010000010";
						 when  154  =>    DADOS_AUDIO <=  "0010101001010000";
						 when  155  =>    DADOS_AUDIO <=  "0010100000011011";
						 when  156  =>    DADOS_AUDIO <=  "0010010111100011";
						 when  157  =>    DADOS_AUDIO <=  "0010001110100111";
						 when  158  =>    DADOS_AUDIO <=  "0010000101101001";
						 when  159  =>    DADOS_AUDIO <=  "0001111100100111";
						 when  160  =>    DADOS_AUDIO <=  "0001110011100011";
						 when  161  =>    DADOS_AUDIO <=  "0001101010011100";
						 when  162  =>    DADOS_AUDIO <=  "0001100001010100";
						 when  163  =>    DADOS_AUDIO <=  "0001011000001001";
						 when  164  =>    DADOS_AUDIO <=  "0001001110111100";
						 when  165  =>    DADOS_AUDIO <=  "0001000101101101";
						 when  166  =>    DADOS_AUDIO <=  "0000111100011101";
						 when  167  =>    DADOS_AUDIO <=  "0000110011001100";
						 when  168  =>    DADOS_AUDIO <=  "0000101001111010";
						 when  169  =>    DADOS_AUDIO <=  "0000100000100111";
						 when  170  =>    DADOS_AUDIO <=  "0000010111010011";
						 when  171  =>    DADOS_AUDIO <=  "0000001101111111";
						 when  172  =>    DADOS_AUDIO <=  "0000000100101010";
						 when  173  =>    DADOS_AUDIO <=  "1111111011010110";
						 when  174  =>    DADOS_AUDIO <=  "1111110010000001";
						 when  175  =>    DADOS_AUDIO <=  "1111101000101101";
						 when  176  =>    DADOS_AUDIO <=  "1111011111011001";
						 when  177  =>    DADOS_AUDIO <=  "1111010110000110";
						 when  178  =>    DADOS_AUDIO <=  "1111001100110100";
						 when  179  =>    DADOS_AUDIO <=  "1111000011100011";
						 when  180  =>    DADOS_AUDIO <=  "1110111010010011";
						 when  181  =>    DADOS_AUDIO <=  "1110110001000100";
						 when  182  =>    DADOS_AUDIO <=  "1110100111110111";
						 when  183  =>    DADOS_AUDIO <=  "1110011110101100";
						 when  184  =>    DADOS_AUDIO <=  "1110010101100100";
						 when  185  =>    DADOS_AUDIO <=  "1110001100011101";
						 when  186  =>    DADOS_AUDIO <=  "1110000011011001";
						 when  187  =>    DADOS_AUDIO <=  "1101111010010111";
						 when  188  =>    DADOS_AUDIO <=  "1101110001011001";
						 when  189  =>    DADOS_AUDIO <=  "1101101000011101";
						 when  190  =>    DADOS_AUDIO <=  "1101011111100101";
						 when  191  =>    DADOS_AUDIO <=  "1101010110110000";
						 when  192  =>    DADOS_AUDIO <=  "1101001101111110";
						 when  193  =>    DADOS_AUDIO <=  "1101000101010001";
						 when  194  =>    DADOS_AUDIO <=  "1100111100100111";
						 when  195  =>    DADOS_AUDIO <=  "1100110100000010";
						 when  196  =>    DADOS_AUDIO <=  "1100101011100001";
						 when  197  =>    DADOS_AUDIO <=  "1100100011000100";
						 when  198  =>    DADOS_AUDIO <=  "1100011010101100";
						 when  199  =>    DADOS_AUDIO <=  "1100010010011001";
						 when  200  =>    DADOS_AUDIO <=  "1100001010001011";
						 when  201  =>    DADOS_AUDIO <=  "1100000010000010";
						 when  202  =>    DADOS_AUDIO <=  "1011111001111110";
						 when  203  =>    DADOS_AUDIO <=  "1011110010000001";
						 when  204  =>    DADOS_AUDIO <=  "1011101010001000";
						 when  205  =>    DADOS_AUDIO <=  "1011100010010110";
						 when  206  =>    DADOS_AUDIO <=  "1011011010101010";
						 when  207  =>    DADOS_AUDIO <=  "1011010011000100";
						 when  208  =>    DADOS_AUDIO <=  "1011001011100100";
						 when  209  =>    DADOS_AUDIO <=  "1011000100001011";
						 when  210  =>    DADOS_AUDIO <=  "1010111100111001";
						 when  211  =>    DADOS_AUDIO <=  "1010110101101110";
						 when  212  =>    DADOS_AUDIO <=  "1010101110101001";
						 when  213  =>    DADOS_AUDIO <=  "1010100111101100";
						 when  214  =>    DADOS_AUDIO <=  "1010100000110110";
						 when  215  =>    DADOS_AUDIO <=  "1010011010000111";
						 when  216  =>    DADOS_AUDIO <=  "1010010011100000";
						 when  217  =>    DADOS_AUDIO <=  "1010001101000001";
						 when  218  =>    DADOS_AUDIO <=  "1010000110101010";
						 when  219  =>    DADOS_AUDIO <=  "1010000000011010";
						 when  220  =>    DADOS_AUDIO <=  "1001111010010011";
						 when  221  =>    DADOS_AUDIO <=  "1001110100010100";
						 when  222  =>    DADOS_AUDIO <=  "1001101110011110";
						 when  223  =>    DADOS_AUDIO <=  "1001101000110000";
						 when  224  =>    DADOS_AUDIO <=  "1001100011001011";
						 when  225  =>    DADOS_AUDIO <=  "1001011101101110";
						 when  226  =>    DADOS_AUDIO <=  "1001011000011010";
						 when  227  =>    DADOS_AUDIO <=  "1001010011010000";
						 when  228  =>    DADOS_AUDIO <=  "1001001110001110";
						 when  229  =>    DADOS_AUDIO <=  "1001001001010110";
						 when  230  =>    DADOS_AUDIO <=  "1001000100100111";
						 when  231  =>    DADOS_AUDIO <=  "1001000000000001";
						 when  232  =>    DADOS_AUDIO <=  "1000111011100101";
						 when  233  =>    DADOS_AUDIO <=  "1000110111010010";
						 when  234  =>    DADOS_AUDIO <=  "1000110011001001";
						 when  235  =>    DADOS_AUDIO <=  "1000101111001010";
						 when  236  =>    DADOS_AUDIO <=  "1000101011010101";
						 when  237  =>    DADOS_AUDIO <=  "1000100111101010";
						 when  238  =>    DADOS_AUDIO <=  "1000100100001001";
						 when  239  =>    DADOS_AUDIO <=  "1000100000110001";
						 when  240  =>    DADOS_AUDIO <=  "1000011101100100";
						 when  241  =>    DADOS_AUDIO <=  "1000011010100010";
						 when  242  =>    DADOS_AUDIO <=  "1000010111101001";
						 when  243  =>    DADOS_AUDIO <=  "1000010100111011";
						 when  244  =>    DADOS_AUDIO <=  "1000010010011000";
						 when  245  =>    DADOS_AUDIO <=  "1000001111111111";
						 when  246  =>    DADOS_AUDIO <=  "1000001101110000";
						 when  247  =>    DADOS_AUDIO <=  "1000001011101100";
						 when  248  =>    DADOS_AUDIO <=  "1000001001110010";
						 when  249  =>    DADOS_AUDIO <=  "1000001000000100";
						 when  250  =>    DADOS_AUDIO <=  "1000000110100000";
						 when  251  =>    DADOS_AUDIO <=  "1000000101000110";
						 when  252  =>    DADOS_AUDIO <=  "1000000011111000";
						 when  253  =>    DADOS_AUDIO <=  "1000000010110100";
						 when  254  =>    DADOS_AUDIO <=  "1000000001111011";
						 when  255  =>    DADOS_AUDIO <=  "1000000001001101";
						 when  256  =>    DADOS_AUDIO <=  "1000000000101010";
						 when  257  =>    DADOS_AUDIO <=  "1000000000010001";
						 when  258  =>    DADOS_AUDIO <=  "1000000000000100";
						 when  259  =>    DADOS_AUDIO <=  "1000000000000001";
						 when  260  =>    DADOS_AUDIO <=  "1000000000001001";
						 when  261  =>    DADOS_AUDIO <=  "1000000000011100";
						 when  262  =>    DADOS_AUDIO <=  "1000000000111010";
						 when  263  =>    DADOS_AUDIO <=  "1000000001100011";
						 when  264  =>    DADOS_AUDIO <=  "1000000010010110";
						 when  265  =>    DADOS_AUDIO <=  "1000000011010101";
						 when  266  =>    DADOS_AUDIO <=  "1000000100011110";
						 when  267  =>    DADOS_AUDIO <=  "1000000101110010";
						 when  268  =>    DADOS_AUDIO <=  "1000000111010000";
						 when  269  =>    DADOS_AUDIO <=  "1000001000111010";
						 when  270  =>    DADOS_AUDIO <=  "1000001010101110";
						 when  271  =>    DADOS_AUDIO <=  "1000001100101101";
						 when  272  =>    DADOS_AUDIO <=  "1000001110110110";
						 when  273  =>    DADOS_AUDIO <=  "1000010001001010";
						 when  274  =>    DADOS_AUDIO <=  "1000010011101000";
						 when  275  =>    DADOS_AUDIO <=  "1000010110010001";
						 when  276  =>    DADOS_AUDIO <=  "1000011001000100";
						 when  277  =>    DADOS_AUDIO <=  "1000011100000010";
						 when  278  =>    DADOS_AUDIO <=  "1000011111001010";
						 when  279  =>    DADOS_AUDIO <=  "1000100010011100";
						 when  280  =>    DADOS_AUDIO <=  "1000100101111000";
						 when  281  =>    DADOS_AUDIO <=  "1000101001011110";
						 when  282  =>    DADOS_AUDIO <=  "1000101101001110";
						 when  283  =>    DADOS_AUDIO <=  "1000110001001001";
						 when  284  =>    DADOS_AUDIO <=  "1000110101001101";
						 when  285  =>    DADOS_AUDIO <=  "1000111001011010";
						 when  286  =>    DADOS_AUDIO <=  "1000111101110010";
						 when  287  =>    DADOS_AUDIO <=  "1001000010010011";
						 when  288  =>    DADOS_AUDIO <=  "1001000110111101";
						 when  289  =>    DADOS_AUDIO <=  "1001001011110001";
						 when  290  =>    DADOS_AUDIO <=  "1001010000101110";
						 when  291  =>    DADOS_AUDIO <=  "1001010101110100";
						 when  292  =>    DADOS_AUDIO <=  "1001011011000011";
						 when  293  =>    DADOS_AUDIO <=  "1001100000011011";
						 when  294  =>    DADOS_AUDIO <=  "1001100101111100";
						 when  295  =>    DADOS_AUDIO <=  "1001101011100110";
						 when  296  =>    DADOS_AUDIO <=  "1001110001011000";
						 when  297  =>    DADOS_AUDIO <=  "1001110111010011";
						 when  298  =>    DADOS_AUDIO <=  "1001111101010110";
						 when  299  =>    DADOS_AUDIO <=  "1010000011100001";
						 when  300  =>    DADOS_AUDIO <=  "1010001001110100";
						 when  301  =>    DADOS_AUDIO <=  "1010010000010000";
						 when  302  =>    DADOS_AUDIO <=  "1010010110110011";
						 when  303  =>    DADOS_AUDIO <=  "1010011101011110";
						 when  304  =>    DADOS_AUDIO <=  "1010100100010000";
						 when  305  =>    DADOS_AUDIO <=  "1010101011001010";
						 when  306  =>    DADOS_AUDIO <=  "1010110010001010";
						 when  307  =>    DADOS_AUDIO <=  "1010111001010010";
						 when  308  =>    DADOS_AUDIO <=  "1011000000100001";
						 when  309  =>    DADOS_AUDIO <=  "1011000111110111";
						 when  310  =>    DADOS_AUDIO <=  "1011001111010011";
						 when  311  =>    DADOS_AUDIO <=  "1011010110110110";
						 when  312  =>    DADOS_AUDIO <=  "1011011110011111";
						 when  313  =>    DADOS_AUDIO <=  "1011100110001110";
						 when  314  =>    DADOS_AUDIO <=  "1011101110000100";
						 when  315  =>    DADOS_AUDIO <=  "1011110101111111";
						 when  316  =>    DADOS_AUDIO <=  "1011111101111111";
						 when  317  =>    DADOS_AUDIO <=  "1100000110000110";
						 when  318  =>    DADOS_AUDIO <=  "1100001110010001";
						 when  319  =>    DADOS_AUDIO <=  "1100010110100010";
						 when  320  =>    DADOS_AUDIO <=  "1100011110110111";
						 when  321  =>    DADOS_AUDIO <=  "1100100111010010";
						 when  322  =>    DADOS_AUDIO <=  "1100101111110001";
						 when  323  =>    DADOS_AUDIO <=  "1100111000010100";
						 when  324  =>    DADOS_AUDIO <=  "1101000000111100";
						 when  325  =>    DADOS_AUDIO <=  "1101001001100111";
						 when  326  =>    DADOS_AUDIO <=  "1101010010010111";
						 when  327  =>    DADOS_AUDIO <=  "1101011011001010";
						 when  328  =>    DADOS_AUDIO <=  "1101100100000001";
						 when  329  =>    DADOS_AUDIO <=  "1101101100111011";
						 when  330  =>    DADOS_AUDIO <=  "1101110101111000";
						 when  331  =>    DADOS_AUDIO <=  "1101111110111000";
						 when  332  =>    DADOS_AUDIO <=  "1110000111111011";
						 when  333  =>    DADOS_AUDIO <=  "1110010001000000";
						 when  334  =>    DADOS_AUDIO <=  "1110011010001000";
						 when  335  =>    DADOS_AUDIO <=  "1110100011010010";
						 when  336  =>    DADOS_AUDIO <=  "1110101100011110";
						 when  337  =>    DADOS_AUDIO <=  "1110110101101011";
						 when  338  =>    DADOS_AUDIO <=  "1110111110111010";
						 when  339  =>    DADOS_AUDIO <=  "1111001000001011";
						 when  340  =>    DADOS_AUDIO <=  "1111010001011101";
						 when  341  =>    DADOS_AUDIO <=  "1111011010110000";
						 when  342  =>    DADOS_AUDIO <=  "1111100100000011";
						 when  343  =>    DADOS_AUDIO <=  "1111101101010111";
						 when  344  =>    DADOS_AUDIO <=  "1111110110101100";
						 when  345  =>    DADOS_AUDIO <=  "0000000000000000";
						 when others =>	DADOS_AUDIO <=  "0000000000000000";
					end case;
				when 3 =>
					n_pontos <= 326;
					reset <= '0';
					case aux_dados is
					    when  0  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  1  =>    DADOS_AUDIO <=  "0000001001111001";
						 when  2  =>    DADOS_AUDIO <=  "0000010011110010";
						 when  3  =>    DADOS_AUDIO <=  "0000011101101011";
						 when  4  =>    DADOS_AUDIO <=  "0000100111100011";
						 when  5  =>    DADOS_AUDIO <=  "0000110001011010";
						 when  6  =>    DADOS_AUDIO <=  "0000111011010000";
						 when  7  =>    DADOS_AUDIO <=  "0001000101000100";
						 when  8  =>    DADOS_AUDIO <=  "0001001110110111";
						 when  9  =>    DADOS_AUDIO <=  "0001011000101000";
						 when  10  =>    DADOS_AUDIO <=  "0001100010010111";
						 when  11  =>    DADOS_AUDIO <=  "0001101100000100";
						 when  12  =>    DADOS_AUDIO <=  "0001110101101101";
						 when  13  =>    DADOS_AUDIO <=  "0001111111010101";
						 when  14  =>    DADOS_AUDIO <=  "0010001000111001";
						 when  15  =>    DADOS_AUDIO <=  "0010010010011001";
						 when  16  =>    DADOS_AUDIO <=  "0010011011110111";
						 when  17  =>    DADOS_AUDIO <=  "0010100101010000";
						 when  18  =>    DADOS_AUDIO <=  "0010101110100110";
						 when  19  =>    DADOS_AUDIO <=  "0010110111110111";
						 when  20  =>    DADOS_AUDIO <=  "0011000001000100";
						 when  21  =>    DADOS_AUDIO <=  "0011001010001101";
						 when  22  =>    DADOS_AUDIO <=  "0011010011010000";
						 when  23  =>    DADOS_AUDIO <=  "0011011100001111";
						 when  24  =>    DADOS_AUDIO <=  "0011100101001000";
						 when  25  =>    DADOS_AUDIO <=  "0011101101111100";
						 when  26  =>    DADOS_AUDIO <=  "0011110110101010";
						 when  27  =>    DADOS_AUDIO <=  "0011111111010010";
						 when  28  =>    DADOS_AUDIO <=  "0100000111110100";
						 when  29  =>    DADOS_AUDIO <=  "0100010000010000";
						 when  30  =>    DADOS_AUDIO <=  "0100011000100101";
						 when  31  =>    DADOS_AUDIO <=  "0100100000110011";
						 when  32  =>    DADOS_AUDIO <=  "0100101000111011";
						 when  33  =>    DADOS_AUDIO <=  "0100110000111011";
						 when  34  =>    DADOS_AUDIO <=  "0100111000110101";
						 when  35  =>    DADOS_AUDIO <=  "0101000000100110";
						 when  36  =>    DADOS_AUDIO <=  "0101001000010000";
						 when  37  =>    DADOS_AUDIO <=  "0101001111110011";
						 when  38  =>    DADOS_AUDIO <=  "0101010111001101";
						 when  39  =>    DADOS_AUDIO <=  "0101011110011111";
						 when  40  =>    DADOS_AUDIO <=  "0101100101101000";
						 when  41  =>    DADOS_AUDIO <=  "0101101100101001";
						 when  42  =>    DADOS_AUDIO <=  "0101110011100010";
						 when  43  =>    DADOS_AUDIO <=  "0101111010010001";
						 when  44  =>    DADOS_AUDIO <=  "0110000000110111";
						 when  45  =>    DADOS_AUDIO <=  "0110000111010101";
						 when  46  =>    DADOS_AUDIO <=  "0110001101101000";
						 when  47  =>    DADOS_AUDIO <=  "0110010011110011";
						 when  48  =>    DADOS_AUDIO <=  "0110011001110011";
						 when  49  =>    DADOS_AUDIO <=  "0110011111101010";
						 when  50  =>    DADOS_AUDIO <=  "0110100101010111";
						 when  51  =>    DADOS_AUDIO <=  "0110101010111010";
						 when  52  =>    DADOS_AUDIO <=  "0110110000010010";
						 when  53  =>    DADOS_AUDIO <=  "0110110101100001";
						 when  54  =>    DADOS_AUDIO <=  "0110111010100100";
						 when  55  =>    DADOS_AUDIO <=  "0110111111011110";
						 when  56  =>    DADOS_AUDIO <=  "0111000100001100";
						 when  57  =>    DADOS_AUDIO <=  "0111001000110000";
						 when  58  =>    DADOS_AUDIO <=  "0111001101001001";
						 when  59  =>    DADOS_AUDIO <=  "0111010001010110";
						 when  60  =>    DADOS_AUDIO <=  "0111010101011001";
						 when  61  =>    DADOS_AUDIO <=  "0111011001010000";
						 when  62  =>    DADOS_AUDIO <=  "0111011100111100";
						 when  63  =>    DADOS_AUDIO <=  "0111100000011101";
						 when  64  =>    DADOS_AUDIO <=  "0111100011110010";
						 when  65  =>    DADOS_AUDIO <=  "0111100110111100";
						 when  66  =>    DADOS_AUDIO <=  "0111101001111010";
						 when  67  =>    DADOS_AUDIO <=  "0111101100101100";
						 when  68  =>    DADOS_AUDIO <=  "0111101111010010";
						 when  69  =>    DADOS_AUDIO <=  "0111110001101101";
						 when  70  =>    DADOS_AUDIO <=  "0111110011111100";
						 when  71  =>    DADOS_AUDIO <=  "0111110101111110";
						 when  72  =>    DADOS_AUDIO <=  "0111110111110101";
						 when  73  =>    DADOS_AUDIO <=  "0111111001100000";
						 when  74  =>    DADOS_AUDIO <=  "0111111010111110";
						 when  75  =>    DADOS_AUDIO <=  "0111111100010001";
						 when  76  =>    DADOS_AUDIO <=  "0111111101010111";
						 when  77  =>    DADOS_AUDIO <=  "0111111110010001";
						 when  78  =>    DADOS_AUDIO <=  "0111111110111111";
						 when  79  =>    DADOS_AUDIO <=  "0111111111100001";
						 when  80  =>    DADOS_AUDIO <=  "0111111111110110";
						 when  81  =>    DADOS_AUDIO <=  "0111111111111111";
						 when  82  =>    DADOS_AUDIO <=  "0111111111111100";
						 when  83  =>    DADOS_AUDIO <=  "0111111111101101";
						 when  84  =>    DADOS_AUDIO <=  "0111111111010001";
						 when  85  =>    DADOS_AUDIO <=  "0111111110101001";
						 when  86  =>    DADOS_AUDIO <=  "0111111101110101";
						 when  87  =>    DADOS_AUDIO <=  "0111111100110101";
						 when  88  =>    DADOS_AUDIO <=  "0111111011101001";
						 when  89  =>    DADOS_AUDIO <=  "0111111010010000";
						 when  90  =>    DADOS_AUDIO <=  "0111111000101100";
						 when  91  =>    DADOS_AUDIO <=  "0111110110111011";
						 when  92  =>    DADOS_AUDIO <=  "0111110100111110";
						 when  93  =>    DADOS_AUDIO <=  "0111110010110110";
						 when  94  =>    DADOS_AUDIO <=  "0111110000100001";
						 when  95  =>    DADOS_AUDIO <=  "0111101110000001";
						 when  96  =>    DADOS_AUDIO <=  "0111101011010100";
						 when  97  =>    DADOS_AUDIO <=  "0111101000011100";
						 when  98  =>    DADOS_AUDIO <=  "0111100101011000";
						 when  99  =>    DADOS_AUDIO <=  "0111100010001001";
						 when  100  =>    DADOS_AUDIO <=  "0111011110101110";
						 when  101  =>    DADOS_AUDIO <=  "0111011011001000";
						 when  102  =>    DADOS_AUDIO <=  "0111010111010110";
						 when  103  =>    DADOS_AUDIO <=  "0111010011011001";
						 when  104  =>    DADOS_AUDIO <=  "0111001111010001";
						 when  105  =>    DADOS_AUDIO <=  "0111001010111110";
						 when  106  =>    DADOS_AUDIO <=  "0111000110011111";
						 when  107  =>    DADOS_AUDIO <=  "0111000001110110";
						 when  108  =>    DADOS_AUDIO <=  "0110111101000010";
						 when  109  =>    DADOS_AUDIO <=  "0110111000000100";
						 when  110  =>    DADOS_AUDIO <=  "0110110010111011";
						 when  111  =>    DADOS_AUDIO <=  "0110101101100111";
						 when  112  =>    DADOS_AUDIO <=  "0110101000001010";
						 when  113  =>    DADOS_AUDIO <=  "0110100010100010";
						 when  114  =>    DADOS_AUDIO <=  "0110011100110000";
						 when  115  =>    DADOS_AUDIO <=  "0110010110110100";
						 when  116  =>    DADOS_AUDIO <=  "0110010000101111";
						 when  117  =>    DADOS_AUDIO <=  "0110001010100000";
						 when  118  =>    DADOS_AUDIO <=  "0110000100000111";
						 when  119  =>    DADOS_AUDIO <=  "0101111101100101";
						 when  120  =>    DADOS_AUDIO <=  "0101110110111010";
						 when  121  =>    DADOS_AUDIO <=  "0101110000000111";
						 when  122  =>    DADOS_AUDIO <=  "0101101001001010";
						 when  123  =>    DADOS_AUDIO <=  "0101100010000101";
						 when  124  =>    DADOS_AUDIO <=  "0101011010110111";
						 when  125  =>    DADOS_AUDIO <=  "0101010011100001";
						 when  126  =>    DADOS_AUDIO <=  "0101001100000010";
						 when  127  =>    DADOS_AUDIO <=  "0101000100011100";
						 when  128  =>    DADOS_AUDIO <=  "0100111100101110";
						 when  129  =>    DADOS_AUDIO <=  "0100110100111001";
						 when  130  =>    DADOS_AUDIO <=  "0100101100111100";
						 when  131  =>    DADOS_AUDIO <=  "0100100100111000";
						 when  132  =>    DADOS_AUDIO <=  "0100011100101101";
						 when  133  =>    DADOS_AUDIO <=  "0100010100011011";
						 when  134  =>    DADOS_AUDIO <=  "0100001100000010";
						 when  135  =>    DADOS_AUDIO <=  "0100000011100100";
						 when  136  =>    DADOS_AUDIO <=  "0011111010111110";
						 when  137  =>    DADOS_AUDIO <=  "0011110010010011";
						 when  138  =>    DADOS_AUDIO <=  "0011101001100010";
						 when  139  =>    DADOS_AUDIO <=  "0011100000101100";
						 when  140  =>    DADOS_AUDIO <=  "0011010111110000";
						 when  141  =>    DADOS_AUDIO <=  "0011001110101111";
						 when  142  =>    DADOS_AUDIO <=  "0011000101101001";
						 when  143  =>    DADOS_AUDIO <=  "0010111100011110";
						 when  144  =>    DADOS_AUDIO <=  "0010110011001111";
						 when  145  =>    DADOS_AUDIO <=  "0010101001111011";
						 when  146  =>    DADOS_AUDIO <=  "0010100000100100";
						 when  147  =>    DADOS_AUDIO <=  "0010010111001000";
						 when  148  =>    DADOS_AUDIO <=  "0010001101101001";
						 when  149  =>    DADOS_AUDIO <=  "0010000100000111";
						 when  150  =>    DADOS_AUDIO <=  "0001111010100001";
						 when  151  =>    DADOS_AUDIO <=  "0001110000111001";
						 when  152  =>    DADOS_AUDIO <=  "0001100111001110";
						 when  153  =>    DADOS_AUDIO <=  "0001011101100000";
						 when  154  =>    DADOS_AUDIO <=  "0001010011110000";
						 when  155  =>    DADOS_AUDIO <=  "0001001001111110";
						 when  156  =>    DADOS_AUDIO <=  "0001000000001010";
						 when  157  =>    DADOS_AUDIO <=  "0000110110010101";
						 when  158  =>    DADOS_AUDIO <=  "0000101100011111";
						 when  159  =>    DADOS_AUDIO <=  "0000100010100111";
						 when  160  =>    DADOS_AUDIO <=  "0000011000101111";
						 when  161  =>    DADOS_AUDIO <=  "0000001110110110";
						 when  162  =>    DADOS_AUDIO <=  "0000000100111100";
						 when  163  =>    DADOS_AUDIO <=  "1111111011000100";
						 when  164  =>    DADOS_AUDIO <=  "1111110001001010";
						 when  165  =>    DADOS_AUDIO <=  "1111100111010001";
						 when  166  =>    DADOS_AUDIO <=  "1111011101011001";
						 when  167  =>    DADOS_AUDIO <=  "1111010011100001";
						 when  168  =>    DADOS_AUDIO <=  "1111001001101011";
						 when  169  =>    DADOS_AUDIO <=  "1110111111110110";
						 when  170  =>    DADOS_AUDIO <=  "1110110110000010";
						 when  171  =>    DADOS_AUDIO <=  "1110101100010000";
						 when  172  =>    DADOS_AUDIO <=  "1110100010100000";
						 when  173  =>    DADOS_AUDIO <=  "1110011000110010";
						 when  174  =>    DADOS_AUDIO <=  "1110001111000111";
						 when  175  =>    DADOS_AUDIO <=  "1110000101011111";
						 when  176  =>    DADOS_AUDIO <=  "1101111011111001";
						 when  177  =>    DADOS_AUDIO <=  "1101110010010111";
						 when  178  =>    DADOS_AUDIO <=  "1101101000111000";
						 when  179  =>    DADOS_AUDIO <=  "1101011111011100";
						 when  180  =>    DADOS_AUDIO <=  "1101010110000101";
						 when  181  =>    DADOS_AUDIO <=  "1101001100110001";
						 when  182  =>    DADOS_AUDIO <=  "1101000011100010";
						 when  183  =>    DADOS_AUDIO <=  "1100111010010111";
						 when  184  =>    DADOS_AUDIO <=  "1100110001010001";
						 when  185  =>    DADOS_AUDIO <=  "1100101000010000";
						 when  186  =>    DADOS_AUDIO <=  "1100011111010100";
						 when  187  =>    DADOS_AUDIO <=  "1100010110011110";
						 when  188  =>    DADOS_AUDIO <=  "1100001101101101";
						 when  189  =>    DADOS_AUDIO <=  "1100000101000010";
						 when  190  =>    DADOS_AUDIO <=  "1011111100011100";
						 when  191  =>    DADOS_AUDIO <=  "1011110011111110";
						 when  192  =>    DADOS_AUDIO <=  "1011101011100101";
						 when  193  =>    DADOS_AUDIO <=  "1011100011010011";
						 when  194  =>    DADOS_AUDIO <=  "1011011011001000";
						 when  195  =>    DADOS_AUDIO <=  "1011010011000100";
						 when  196  =>    DADOS_AUDIO <=  "1011001011000111";
						 when  197  =>    DADOS_AUDIO <=  "1011000011010010";
						 when  198  =>    DADOS_AUDIO <=  "1010111011100100";
						 when  199  =>    DADOS_AUDIO <=  "1010110011111110";
						 when  200  =>    DADOS_AUDIO <=  "1010101100011111";
						 when  201  =>    DADOS_AUDIO <=  "1010100101001001";
						 when  202  =>    DADOS_AUDIO <=  "1010011101111011";
						 when  203  =>    DADOS_AUDIO <=  "1010010110110110";
						 when  204  =>    DADOS_AUDIO <=  "1010001111111001";
						 when  205  =>    DADOS_AUDIO <=  "1010001001000110";
						 when  206  =>    DADOS_AUDIO <=  "1010000010011011";
						 when  207  =>    DADOS_AUDIO <=  "1001111011111001";
						 when  208  =>    DADOS_AUDIO <=  "1001110101100000";
						 when  209  =>    DADOS_AUDIO <=  "1001101111010001";
						 when  210  =>    DADOS_AUDIO <=  "1001101001001100";
						 when  211  =>    DADOS_AUDIO <=  "1001100011010000";
						 when  212  =>    DADOS_AUDIO <=  "1001011101011110";
						 when  213  =>    DADOS_AUDIO <=  "1001010111110110";
						 when  214  =>    DADOS_AUDIO <=  "1001010010011001";
						 when  215  =>    DADOS_AUDIO <=  "1001001101000101";
						 when  216  =>    DADOS_AUDIO <=  "1001000111111100";
						 when  217  =>    DADOS_AUDIO <=  "1001000010111110";
						 when  218  =>    DADOS_AUDIO <=  "1000111110001010";
						 when  219  =>    DADOS_AUDIO <=  "1000111001100001";
						 when  220  =>    DADOS_AUDIO <=  "1000110101000010";
						 when  221  =>    DADOS_AUDIO <=  "1000110000101111";
						 when  222  =>    DADOS_AUDIO <=  "1000101100100111";
						 when  223  =>    DADOS_AUDIO <=  "1000101000101010";
						 when  224  =>    DADOS_AUDIO <=  "1000100100111000";
						 when  225  =>    DADOS_AUDIO <=  "1000100001010010";
						 when  226  =>    DADOS_AUDIO <=  "1000011101110111";
						 when  227  =>    DADOS_AUDIO <=  "1000011010101000";
						 when  228  =>    DADOS_AUDIO <=  "1000010111100100";
						 when  229  =>    DADOS_AUDIO <=  "1000010100101100";
						 when  230  =>    DADOS_AUDIO <=  "1000010001111111";
						 when  231  =>    DADOS_AUDIO <=  "1000001111011111";
						 when  232  =>    DADOS_AUDIO <=  "1000001101001010";
						 when  233  =>    DADOS_AUDIO <=  "1000001011000010";
						 when  234  =>    DADOS_AUDIO <=  "1000001001000101";
						 when  235  =>    DADOS_AUDIO <=  "1000000111010100";
						 when  236  =>    DADOS_AUDIO <=  "1000000101110000";
						 when  237  =>    DADOS_AUDIO <=  "1000000100010111";
						 when  238  =>    DADOS_AUDIO <=  "1000000011001011";
						 when  239  =>    DADOS_AUDIO <=  "1000000010001011";
						 when  240  =>    DADOS_AUDIO <=  "1000000001010111";
						 when  241  =>    DADOS_AUDIO <=  "1000000000101111";
						 when  242  =>    DADOS_AUDIO <=  "1000000000010011";
						 when  243  =>    DADOS_AUDIO <=  "1000000000000100";
						 when  244  =>    DADOS_AUDIO <=  "1000000000000001";
						 when  245  =>    DADOS_AUDIO <=  "1000000000001010";
						 when  246  =>    DADOS_AUDIO <=  "1000000000011111";
						 when  247  =>    DADOS_AUDIO <=  "1000000001000001";
						 when  248  =>    DADOS_AUDIO <=  "1000000001101111";
						 when  249  =>    DADOS_AUDIO <=  "1000000010101001";
						 when  250  =>    DADOS_AUDIO <=  "1000000011101111";
						 when  251  =>    DADOS_AUDIO <=  "1000000101000010";
						 when  252  =>    DADOS_AUDIO <=  "1000000110100000";
						 when  253  =>    DADOS_AUDIO <=  "1000001000001011";
						 when  254  =>    DADOS_AUDIO <=  "1000001010000010";
						 when  255  =>    DADOS_AUDIO <=  "1000001100000100";
						 when  256  =>    DADOS_AUDIO <=  "1000001110010011";
						 when  257  =>    DADOS_AUDIO <=  "1000010000101110";
						 when  258  =>    DADOS_AUDIO <=  "1000010011010100";
						 when  259  =>    DADOS_AUDIO <=  "1000010110000110";
						 when  260  =>    DADOS_AUDIO <=  "1000011001000100";
						 when  261  =>    DADOS_AUDIO <=  "1000011100001110";
						 when  262  =>    DADOS_AUDIO <=  "1000011111100011";
						 when  263  =>    DADOS_AUDIO <=  "1000100011000100";
						 when  264  =>    DADOS_AUDIO <=  "1000100110110000";
						 when  265  =>    DADOS_AUDIO <=  "1000101010100111";
						 when  266  =>    DADOS_AUDIO <=  "1000101110101010";
						 when  267  =>    DADOS_AUDIO <=  "1000110010110111";
						 when  268  =>    DADOS_AUDIO <=  "1000110111010000";
						 when  269  =>    DADOS_AUDIO <=  "1000111011110100";
						 when  270  =>    DADOS_AUDIO <=  "1001000000100010";
						 when  271  =>    DADOS_AUDIO <=  "1001000101011100";
						 when  272  =>    DADOS_AUDIO <=  "1001001010011111";
						 when  273  =>    DADOS_AUDIO <=  "1001001111101110";
						 when  274  =>    DADOS_AUDIO <=  "1001010101000110";
						 when  275  =>    DADOS_AUDIO <=  "1001011010101001";
						 when  276  =>    DADOS_AUDIO <=  "1001100000010110";
						 when  277  =>    DADOS_AUDIO <=  "1001100110001101";
						 when  278  =>    DADOS_AUDIO <=  "1001101100001101";
						 when  279  =>    DADOS_AUDIO <=  "1001110010011000";
						 when  280  =>    DADOS_AUDIO <=  "1001111000101011";
						 when  281  =>    DADOS_AUDIO <=  "1001111111001001";
						 when  282  =>    DADOS_AUDIO <=  "1010000101101111";
						 when  283  =>    DADOS_AUDIO <=  "1010001100011110";
						 when  284  =>    DADOS_AUDIO <=  "1010010011010111";
						 when  285  =>    DADOS_AUDIO <=  "1010011010011000";
						 when  286  =>    DADOS_AUDIO <=  "1010100001100001";
						 when  287  =>    DADOS_AUDIO <=  "1010101000110011";
						 when  288  =>    DADOS_AUDIO <=  "1010110000001101";
						 when  289  =>    DADOS_AUDIO <=  "1010110111110000";
						 when  290  =>    DADOS_AUDIO <=  "1010111111011010";
						 when  291  =>    DADOS_AUDIO <=  "1011000111001011";
						 when  292  =>    DADOS_AUDIO <=  "1011001111000101";
						 when  293  =>    DADOS_AUDIO <=  "1011010111000101";
						 when  294  =>    DADOS_AUDIO <=  "1011011111001101";
						 when  295  =>    DADOS_AUDIO <=  "1011100111011011";
						 when  296  =>    DADOS_AUDIO <=  "1011101111110000";
						 when  297  =>    DADOS_AUDIO <=  "1011111000001100";
						 when  298  =>    DADOS_AUDIO <=  "1100000000101110";
						 when  299  =>    DADOS_AUDIO <=  "1100001001010110";
						 when  300  =>    DADOS_AUDIO <=  "1100010010000100";
						 when  301  =>    DADOS_AUDIO <=  "1100011010111000";
						 when  302  =>    DADOS_AUDIO <=  "1100100011110001";
						 when  303  =>    DADOS_AUDIO <=  "1100101100110000";
						 when  304  =>    DADOS_AUDIO <=  "1100110101110011";
						 when  305  =>    DADOS_AUDIO <=  "1100111110111100";
						 when  306  =>    DADOS_AUDIO <=  "1101001000001001";
						 when  307  =>    DADOS_AUDIO <=  "1101010001011010";
						 when  308  =>    DADOS_AUDIO <=  "1101011010110000";
						 when  309  =>    DADOS_AUDIO <=  "1101100100001001";
						 when  310  =>    DADOS_AUDIO <=  "1101101101100111";
						 when  311  =>    DADOS_AUDIO <=  "1101110111000111";
						 when  312  =>    DADOS_AUDIO <=  "1110000000101011";
						 when  313  =>    DADOS_AUDIO <=  "1110001010010011";
						 when  314  =>    DADOS_AUDIO <=  "1110010011111100";
						 when  315  =>    DADOS_AUDIO <=  "1110011101101001";
						 when  316  =>    DADOS_AUDIO <=  "1110100111011000";
						 when  317  =>    DADOS_AUDIO <=  "1110110001001001";
						 when  318  =>    DADOS_AUDIO <=  "1110111010111100";
						 when  319  =>    DADOS_AUDIO <=  "1111000100110000";
						 when  320  =>    DADOS_AUDIO <=  "1111001110100110";
						 when  321  =>    DADOS_AUDIO <=  "1111011000011101";
						 when  322  =>    DADOS_AUDIO <=  "1111100010010101";
						 when  323  =>    DADOS_AUDIO <=  "1111101100001110";
						 when  324  =>    DADOS_AUDIO <=  "1111110110000111";
						 when  325  =>    DADOS_AUDIO <=  "0000000000000000";
						 when others =>	DADOS_AUDIO <=  "0000000000000000";
					end case;
				when 4 =>
					n_pontos <= 308;
					reset <= '0';
					case aux_dados is
					    when  0  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  1  =>    DADOS_AUDIO <=  "0000001010011110";
						 when  2  =>    DADOS_AUDIO <=  "0000010100111100";
						 when  3  =>    DADOS_AUDIO <=  "0000011111011010";
						 when  4  =>    DADOS_AUDIO <=  "0000101001110111";
						 when  5  =>    DADOS_AUDIO <=  "0000110100010011";
						 when  6  =>    DADOS_AUDIO <=  "0000111110101101";
						 when  7  =>    DADOS_AUDIO <=  "0001001001000110";
						 when  8  =>    DADOS_AUDIO <=  "0001010011011101";
						 when  9  =>    DADOS_AUDIO <=  "0001011101110001";
						 when  10  =>    DADOS_AUDIO <=  "0001101000000011";
						 when  11  =>    DADOS_AUDIO <=  "0001110010010010";
						 when  12  =>    DADOS_AUDIO <=  "0001111100011111";
						 when  13  =>    DADOS_AUDIO <=  "0010000110100111";
						 when  14  =>    DADOS_AUDIO <=  "0010010000101101";
						 when  15  =>    DADOS_AUDIO <=  "0010011010101110";
						 when  16  =>    DADOS_AUDIO <=  "0010100100101011";
						 when  17  =>    DADOS_AUDIO <=  "0010101110100100";
						 when  18  =>    DADOS_AUDIO <=  "0010111000011000";
						 when  19  =>    DADOS_AUDIO <=  "0011000010000111";
						 when  20  =>    DADOS_AUDIO <=  "0011001011110001";
						 when  21  =>    DADOS_AUDIO <=  "0011010101010101";
						 when  22  =>    DADOS_AUDIO <=  "0011011110110100";
						 when  23  =>    DADOS_AUDIO <=  "0011101000001101";
						 when  24  =>    DADOS_AUDIO <=  "0011110001011111";
						 when  25  =>    DADOS_AUDIO <=  "0011111010101100";
						 when  26  =>    DADOS_AUDIO <=  "0100000011110001";
						 when  27  =>    DADOS_AUDIO <=  "0100001100101111";
						 when  28  =>    DADOS_AUDIO <=  "0100010101100110";
						 when  29  =>    DADOS_AUDIO <=  "0100011110010110";
						 when  30  =>    DADOS_AUDIO <=  "0100100110111110";
						 when  31  =>    DADOS_AUDIO <=  "0100101111011110";
						 when  32  =>    DADOS_AUDIO <=  "0100110111110110";
						 when  33  =>    DADOS_AUDIO <=  "0101000000000110";
						 when  34  =>    DADOS_AUDIO <=  "0101001000001101";
						 when  35  =>    DADOS_AUDIO <=  "0101010000001100";
						 when  36  =>    DADOS_AUDIO <=  "0101011000000001";
						 when  37  =>    DADOS_AUDIO <=  "0101011111101101";
						 when  38  =>    DADOS_AUDIO <=  "0101100111001111";
						 when  39  =>    DADOS_AUDIO <=  "0101101110101000";
						 when  40  =>    DADOS_AUDIO <=  "0101110101111000";
						 when  41  =>    DADOS_AUDIO <=  "0101111100111101";
						 when  42  =>    DADOS_AUDIO <=  "0110000011111000";
						 when  43  =>    DADOS_AUDIO <=  "0110001010101000";
						 when  44  =>    DADOS_AUDIO <=  "0110010001001110";
						 when  45  =>    DADOS_AUDIO <=  "0110010111101001";
						 when  46  =>    DADOS_AUDIO <=  "0110011101111010";
						 when  47  =>    DADOS_AUDIO <=  "0110100011111111";
						 when  48  =>    DADOS_AUDIO <=  "0110101001111001";
						 when  49  =>    DADOS_AUDIO <=  "0110101111100111";
						 when  50  =>    DADOS_AUDIO <=  "0110110101001010";
						 when  51  =>    DADOS_AUDIO <=  "0110111010100001";
						 when  52  =>    DADOS_AUDIO <=  "0110111111101101";
						 when  53  =>    DADOS_AUDIO <=  "0111000100101100";
						 when  54  =>    DADOS_AUDIO <=  "0111001001011111";
						 when  55  =>    DADOS_AUDIO <=  "0111001110000110";
						 when  56  =>    DADOS_AUDIO <=  "0111010010100001";
						 when  57  =>    DADOS_AUDIO <=  "0111010110101111";
						 when  58  =>    DADOS_AUDIO <=  "0111011010110000";
						 when  59  =>    DADOS_AUDIO <=  "0111011110100101";
						 when  60  =>    DADOS_AUDIO <=  "0111100010001101";
						 when  61  =>    DADOS_AUDIO <=  "0111100101101000";
						 when  62  =>    DADOS_AUDIO <=  "0111101000110110";
						 when  63  =>    DADOS_AUDIO <=  "0111101011110111";
						 when  64  =>    DADOS_AUDIO <=  "0111101110101010";
						 when  65  =>    DADOS_AUDIO <=  "0111110001010001";
						 when  66  =>    DADOS_AUDIO <=  "0111110011101010";
						 when  67  =>    DADOS_AUDIO <=  "0111110101110101";
						 when  68  =>    DADOS_AUDIO <=  "0111110111110011";
						 when  69  =>    DADOS_AUDIO <=  "0111111001100100";
						 when  70  =>    DADOS_AUDIO <=  "0111111011000111";
						 when  71  =>    DADOS_AUDIO <=  "0111111100011101";
						 when  72  =>    DADOS_AUDIO <=  "0111111101100101";
						 when  73  =>    DADOS_AUDIO <=  "0111111110011111";
						 when  74  =>    DADOS_AUDIO <=  "0111111111001100";
						 when  75  =>    DADOS_AUDIO <=  "0111111111101010";
						 when  76  =>    DADOS_AUDIO <=  "0111111111111100";
						 when  77  =>    DADOS_AUDIO <=  "0111111111111111";
						 when  78  =>    DADOS_AUDIO <=  "0111111111110101";
						 when  79  =>    DADOS_AUDIO <=  "0111111111011101";
						 when  80  =>    DADOS_AUDIO <=  "0111111110110111";
						 when  81  =>    DADOS_AUDIO <=  "0111111110000100";
						 when  82  =>    DADOS_AUDIO <=  "0111111101000011";
						 when  83  =>    DADOS_AUDIO <=  "0111111011110100";
						 when  84  =>    DADOS_AUDIO <=  "0111111010010111";
						 when  85  =>    DADOS_AUDIO <=  "0111111000101110";
						 when  86  =>    DADOS_AUDIO <=  "0111110110110110";
						 when  87  =>    DADOS_AUDIO <=  "0111110100110001";
						 when  88  =>    DADOS_AUDIO <=  "0111110010011111";
						 when  89  =>    DADOS_AUDIO <=  "0111101111111111";
						 when  90  =>    DADOS_AUDIO <=  "0111101101010010";
						 when  91  =>    DADOS_AUDIO <=  "0111101010011000";
						 when  92  =>    DADOS_AUDIO <=  "0111100111010000";
						 when  93  =>    DADOS_AUDIO <=  "0111100011111100";
						 when  94  =>    DADOS_AUDIO <=  "0111100000011011";
						 when  95  =>    DADOS_AUDIO <=  "0111011100101100";
						 when  96  =>    DADOS_AUDIO <=  "0111011000110001";
						 when  97  =>    DADOS_AUDIO <=  "0111010100101001";
						 when  98  =>    DADOS_AUDIO <=  "0111010000010101";
						 when  99  =>    DADOS_AUDIO <=  "0111001011110100";
						 when  100  =>    DADOS_AUDIO <=  "0111000111000111";
						 when  101  =>    DADOS_AUDIO <=  "0111000010001110";
						 when  102  =>    DADOS_AUDIO <=  "0110111101001001";
						 when  103  =>    DADOS_AUDIO <=  "0110110111110111";
						 when  104  =>    DADOS_AUDIO <=  "0110110010011010";
						 when  105  =>    DADOS_AUDIO <=  "0110101100110001";
						 when  106  =>    DADOS_AUDIO <=  "0110100110111101";
						 when  107  =>    DADOS_AUDIO <=  "0110100000111110";
						 when  108  =>    DADOS_AUDIO <=  "0110011010110011";
						 when  109  =>    DADOS_AUDIO <=  "0110010100011101";
						 when  110  =>    DADOS_AUDIO <=  "0110001101111101";
						 when  111  =>    DADOS_AUDIO <=  "0110000111010001";
						 when  112  =>    DADOS_AUDIO <=  "0110000000011100";
						 when  113  =>    DADOS_AUDIO <=  "0101111001011011";
						 when  114  =>    DADOS_AUDIO <=  "0101110010010001";
						 when  115  =>    DADOS_AUDIO <=  "0101101010111101";
						 when  116  =>    DADOS_AUDIO <=  "0101100011011111";
						 when  117  =>    DADOS_AUDIO <=  "0101011011111000";
						 when  118  =>    DADOS_AUDIO <=  "0101010100000111";
						 when  119  =>    DADOS_AUDIO <=  "0101001100001101";
						 when  120  =>    DADOS_AUDIO <=  "0101000100001011";
						 when  121  =>    DADOS_AUDIO <=  "0100111011111111";
						 when  122  =>    DADOS_AUDIO <=  "0100110011101011";
						 when  123  =>    DADOS_AUDIO <=  "0100101011001111";
						 when  124  =>    DADOS_AUDIO <=  "0100100010101011";
						 when  125  =>    DADOS_AUDIO <=  "0100011001111111";
						 when  126  =>    DADOS_AUDIO <=  "0100010001001100";
						 when  127  =>    DADOS_AUDIO <=  "0100001000010001";
						 when  128  =>    DADOS_AUDIO <=  "0011111111001111";
						 when  129  =>    DADOS_AUDIO <=  "0011110110000110";
						 when  130  =>    DADOS_AUDIO <=  "0011101100110111";
						 when  131  =>    DADOS_AUDIO <=  "0011100011100001";
						 when  132  =>    DADOS_AUDIO <=  "0011011010000110";
						 when  133  =>    DADOS_AUDIO <=  "0011010000100100";
						 when  134  =>    DADOS_AUDIO <=  "0011000110111101";
						 when  135  =>    DADOS_AUDIO <=  "0010111101010000";
						 when  136  =>    DADOS_AUDIO <=  "0010110011011110";
						 when  137  =>    DADOS_AUDIO <=  "0010101001101000";
						 when  138  =>    DADOS_AUDIO <=  "0010011111101101";
						 when  139  =>    DADOS_AUDIO <=  "0010010101101110";
						 when  140  =>    DADOS_AUDIO <=  "0010001011101010";
						 when  141  =>    DADOS_AUDIO <=  "0010000001100011";
						 when  142  =>    DADOS_AUDIO <=  "0001110111011001";
						 when  143  =>    DADOS_AUDIO <=  "0001101101001011";
						 when  144  =>    DADOS_AUDIO <=  "0001100010111011";
						 when  145  =>    DADOS_AUDIO <=  "0001011000100111";
						 when  146  =>    DADOS_AUDIO <=  "0001001110010010";
						 when  147  =>    DADOS_AUDIO <=  "0001000011111010";
						 when  148  =>    DADOS_AUDIO <=  "0000111001100000";
						 when  149  =>    DADOS_AUDIO <=  "0000101111000101";
						 when  150  =>    DADOS_AUDIO <=  "0000100100101001";
						 when  151  =>    DADOS_AUDIO <=  "0000011010001011";
						 when  152  =>    DADOS_AUDIO <=  "0000001111101101";
						 when  153  =>    DADOS_AUDIO <=  "0000000101001111";
						 when  154  =>    DADOS_AUDIO <=  "1111111010110001";
						 when  155  =>    DADOS_AUDIO <=  "1111110000010011";
						 when  156  =>    DADOS_AUDIO <=  "1111100101110101";
						 when  157  =>    DADOS_AUDIO <=  "1111011011010111";
						 when  158  =>    DADOS_AUDIO <=  "1111010000111011";
						 when  159  =>    DADOS_AUDIO <=  "1111000110100000";
						 when  160  =>    DADOS_AUDIO <=  "1110111100000110";
						 when  161  =>    DADOS_AUDIO <=  "1110110001101110";
						 when  162  =>    DADOS_AUDIO <=  "1110100111011001";
						 when  163  =>    DADOS_AUDIO <=  "1110011101000101";
						 when  164  =>    DADOS_AUDIO <=  "1110010010110101";
						 when  165  =>    DADOS_AUDIO <=  "1110001000100111";
						 when  166  =>    DADOS_AUDIO <=  "1101111110011101";
						 when  167  =>    DADOS_AUDIO <=  "1101110100010110";
						 when  168  =>    DADOS_AUDIO <=  "1101101010010010";
						 when  169  =>    DADOS_AUDIO <=  "1101100000010011";
						 when  170  =>    DADOS_AUDIO <=  "1101010110011000";
						 when  171  =>    DADOS_AUDIO <=  "1101001100100010";
						 when  172  =>    DADOS_AUDIO <=  "1101000010110000";
						 when  173  =>    DADOS_AUDIO <=  "1100111001000011";
						 when  174  =>    DADOS_AUDIO <=  "1100101111011100";
						 when  175  =>    DADOS_AUDIO <=  "1100100101111010";
						 when  176  =>    DADOS_AUDIO <=  "1100011100011111";
						 when  177  =>    DADOS_AUDIO <=  "1100010011001001";
						 when  178  =>    DADOS_AUDIO <=  "1100001001111010";
						 when  179  =>    DADOS_AUDIO <=  "1100000000110001";
						 when  180  =>    DADOS_AUDIO <=  "1011110111101111";
						 when  181  =>    DADOS_AUDIO <=  "1011101110110100";
						 when  182  =>    DADOS_AUDIO <=  "1011100110000001";
						 when  183  =>    DADOS_AUDIO <=  "1011011101010101";
						 when  184  =>    DADOS_AUDIO <=  "1011010100110001";
						 when  185  =>    DADOS_AUDIO <=  "1011001100010101";
						 when  186  =>    DADOS_AUDIO <=  "1011000100000001";
						 when  187  =>    DADOS_AUDIO <=  "1010111011110101";
						 when  188  =>    DADOS_AUDIO <=  "1010110011110011";
						 when  189  =>    DADOS_AUDIO <=  "1010101011111001";
						 when  190  =>    DADOS_AUDIO <=  "1010100100001000";
						 when  191  =>    DADOS_AUDIO <=  "1010011100100001";
						 when  192  =>    DADOS_AUDIO <=  "1010010101000011";
						 when  193  =>    DADOS_AUDIO <=  "1010001101101111";
						 when  194  =>    DADOS_AUDIO <=  "1010000110100101";
						 when  195  =>    DADOS_AUDIO <=  "1001111111100100";
						 when  196  =>    DADOS_AUDIO <=  "1001111000101111";
						 when  197  =>    DADOS_AUDIO <=  "1001110010000011";
						 when  198  =>    DADOS_AUDIO <=  "1001101011100011";
						 when  199  =>    DADOS_AUDIO <=  "1001100101001101";
						 when  200  =>    DADOS_AUDIO <=  "1001011111000010";
						 when  201  =>    DADOS_AUDIO <=  "1001011001000011";
						 when  202  =>    DADOS_AUDIO <=  "1001010011001111";
						 when  203  =>    DADOS_AUDIO <=  "1001001101100110";
						 when  204  =>    DADOS_AUDIO <=  "1001001000001001";
						 when  205  =>    DADOS_AUDIO <=  "1001000010110111";
						 when  206  =>    DADOS_AUDIO <=  "1000111101110010";
						 when  207  =>    DADOS_AUDIO <=  "1000111000111001";
						 when  208  =>    DADOS_AUDIO <=  "1000110100001100";
						 when  209  =>    DADOS_AUDIO <=  "1000101111101011";
						 when  210  =>    DADOS_AUDIO <=  "1000101011010111";
						 when  211  =>    DADOS_AUDIO <=  "1000100111001111";
						 when  212  =>    DADOS_AUDIO <=  "1000100011010100";
						 when  213  =>    DADOS_AUDIO <=  "1000011111100101";
						 when  214  =>    DADOS_AUDIO <=  "1000011100000100";
						 when  215  =>    DADOS_AUDIO <=  "1000011000110000";
						 when  216  =>    DADOS_AUDIO <=  "1000010101101000";
						 when  217  =>    DADOS_AUDIO <=  "1000010010101110";
						 when  218  =>    DADOS_AUDIO <=  "1000010000000001";
						 when  219  =>    DADOS_AUDIO <=  "1000001101100001";
						 when  220  =>    DADOS_AUDIO <=  "1000001011001111";
						 when  221  =>    DADOS_AUDIO <=  "1000001001001010";
						 when  222  =>    DADOS_AUDIO <=  "1000000111010010";
						 when  223  =>    DADOS_AUDIO <=  "1000000101101001";
						 when  224  =>    DADOS_AUDIO <=  "1000000100001100";
						 when  225  =>    DADOS_AUDIO <=  "1000000010111101";
						 when  226  =>    DADOS_AUDIO <=  "1000000001111100";
						 when  227  =>    DADOS_AUDIO <=  "1000000001001001";
						 when  228  =>    DADOS_AUDIO <=  "1000000000100011";
						 when  229  =>    DADOS_AUDIO <=  "1000000000001011";
						 when  230  =>    DADOS_AUDIO <=  "1000000000000001";
						 when  231  =>    DADOS_AUDIO <=  "1000000000000100";
						 when  232  =>    DADOS_AUDIO <=  "1000000000010110";
						 when  233  =>    DADOS_AUDIO <=  "1000000000110100";
						 when  234  =>    DADOS_AUDIO <=  "1000000001100001";
						 when  235  =>    DADOS_AUDIO <=  "1000000010011011";
						 when  236  =>    DADOS_AUDIO <=  "1000000011100011";
						 when  237  =>    DADOS_AUDIO <=  "1000000100111001";
						 when  238  =>    DADOS_AUDIO <=  "1000000110011100";
						 when  239  =>    DADOS_AUDIO <=  "1000001000001101";
						 when  240  =>    DADOS_AUDIO <=  "1000001010001011";
						 when  241  =>    DADOS_AUDIO <=  "1000001100010110";
						 when  242  =>    DADOS_AUDIO <=  "1000001110101111";
						 when  243  =>    DADOS_AUDIO <=  "1000010001010110";
						 when  244  =>    DADOS_AUDIO <=  "1000010100001001";
						 when  245  =>    DADOS_AUDIO <=  "1000010111001010";
						 when  246  =>    DADOS_AUDIO <=  "1000011010011000";
						 when  247  =>    DADOS_AUDIO <=  "1000011101110011";
						 when  248  =>    DADOS_AUDIO <=  "1000100001011011";
						 when  249  =>    DADOS_AUDIO <=  "1000100101010000";
						 when  250  =>    DADOS_AUDIO <=  "1000101001010001";
						 when  251  =>    DADOS_AUDIO <=  "1000101101011111";
						 when  252  =>    DADOS_AUDIO <=  "1000110001111010";
						 when  253  =>    DADOS_AUDIO <=  "1000110110100001";
						 when  254  =>    DADOS_AUDIO <=  "1000111011010100";
						 when  255  =>    DADOS_AUDIO <=  "1001000000010011";
						 when  256  =>    DADOS_AUDIO <=  "1001000101011111";
						 when  257  =>    DADOS_AUDIO <=  "1001001010110110";
						 when  258  =>    DADOS_AUDIO <=  "1001010000011001";
						 when  259  =>    DADOS_AUDIO <=  "1001010110000111";
						 when  260  =>    DADOS_AUDIO <=  "1001011100000001";
						 when  261  =>    DADOS_AUDIO <=  "1001100010000110";
						 when  262  =>    DADOS_AUDIO <=  "1001101000010111";
						 when  263  =>    DADOS_AUDIO <=  "1001101110110010";
						 when  264  =>    DADOS_AUDIO <=  "1001110101011000";
						 when  265  =>    DADOS_AUDIO <=  "1001111100001000";
						 when  266  =>    DADOS_AUDIO <=  "1010000011000011";
						 when  267  =>    DADOS_AUDIO <=  "1010001010001000";
						 when  268  =>    DADOS_AUDIO <=  "1010010001011000";
						 when  269  =>    DADOS_AUDIO <=  "1010011000110001";
						 when  270  =>    DADOS_AUDIO <=  "1010100000010011";
						 when  271  =>    DADOS_AUDIO <=  "1010100111111111";
						 when  272  =>    DADOS_AUDIO <=  "1010101111110100";
						 when  273  =>    DADOS_AUDIO <=  "1010110111110011";
						 when  274  =>    DADOS_AUDIO <=  "1010111111111010";
						 when  275  =>    DADOS_AUDIO <=  "1011001000001010";
						 when  276  =>    DADOS_AUDIO <=  "1011010000100010";
						 when  277  =>    DADOS_AUDIO <=  "1011011001000010";
						 when  278  =>    DADOS_AUDIO <=  "1011100001101010";
						 when  279  =>    DADOS_AUDIO <=  "1011101010011010";
						 when  280  =>    DADOS_AUDIO <=  "1011110011010001";
						 when  281  =>    DADOS_AUDIO <=  "1011111100001111";
						 when  282  =>    DADOS_AUDIO <=  "1100000101010100";
						 when  283  =>    DADOS_AUDIO <=  "1100001110100001";
						 when  284  =>    DADOS_AUDIO <=  "1100010111110011";
						 when  285  =>    DADOS_AUDIO <=  "1100100001001100";
						 when  286  =>    DADOS_AUDIO <=  "1100101010101011";
						 when  287  =>    DADOS_AUDIO <=  "1100110100001111";
						 when  288  =>    DADOS_AUDIO <=  "1100111101111001";
						 when  289  =>    DADOS_AUDIO <=  "1101000111101000";
						 when  290  =>    DADOS_AUDIO <=  "1101010001011100";
						 when  291  =>    DADOS_AUDIO <=  "1101011011010101";
						 when  292  =>    DADOS_AUDIO <=  "1101100101010010";
						 when  293  =>    DADOS_AUDIO <=  "1101101111010011";
						 when  294  =>    DADOS_AUDIO <=  "1101111001011001";
						 when  295  =>    DADOS_AUDIO <=  "1110000011100001";
						 when  296  =>    DADOS_AUDIO <=  "1110001101101110";
						 when  297  =>    DADOS_AUDIO <=  "1110010111111101";
						 when  298  =>    DADOS_AUDIO <=  "1110100010001111";
						 when  299  =>    DADOS_AUDIO <=  "1110101100100011";
						 when  300  =>    DADOS_AUDIO <=  "1110110110111010";
						 when  301  =>    DADOS_AUDIO <=  "1111000001010011";
						 when  302  =>    DADOS_AUDIO <=  "1111001011101101";
						 when  303  =>    DADOS_AUDIO <=  "1111010110001001";
						 when  304  =>    DADOS_AUDIO <=  "1111100000100110";
						 when  305  =>    DADOS_AUDIO <=  "1111101011000100";
						 when  306  =>    DADOS_AUDIO <=  "1111110101100010";
						 when  307  =>    DADOS_AUDIO <=  "0000000000000000";
						 when others =>	DADOS_AUDIO <=  "0000000000000000";
					end case;
				when 5 =>
					n_pontos <= 290;
					reset <= '0';
					case aux_dados is
					    when  0  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  1  =>    DADOS_AUDIO <=  "0000001011001000";
						 when  2  =>    DADOS_AUDIO <=  "0000010110010000";
						 when  3  =>    DADOS_AUDIO <=  "0000100001010111";
						 when  4  =>    DADOS_AUDIO <=  "0000101100011110";
						 when  5  =>    DADOS_AUDIO <=  "0000110111100011";
						 when  6  =>    DADOS_AUDIO <=  "0001000010100110";
						 when  7  =>    DADOS_AUDIO <=  "0001001101100111";
						 when  8  =>    DADOS_AUDIO <=  "0001011000100110";
						 when  9  =>    DADOS_AUDIO <=  "0001100011100010";
						 when  10  =>    DADOS_AUDIO <=  "0001101110011100";
						 when  11  =>    DADOS_AUDIO <=  "0001111001010010";
						 when  12  =>    DADOS_AUDIO <=  "0010000100000100";
						 when  13  =>    DADOS_AUDIO <=  "0010001110110010";
						 when  14  =>    DADOS_AUDIO <=  "0010011001011100";
						 when  15  =>    DADOS_AUDIO <=  "0010100100000001";
						 when  16  =>    DADOS_AUDIO <=  "0010101110100010";
						 when  17  =>    DADOS_AUDIO <=  "0010111000111101";
						 when  18  =>    DADOS_AUDIO <=  "0011000011010010";
						 when  19  =>    DADOS_AUDIO <=  "0011001101100010";
						 when  20  =>    DADOS_AUDIO <=  "0011010111101011";
						 when  21  =>    DADOS_AUDIO <=  "0011100001101110";
						 when  22  =>    DADOS_AUDIO <=  "0011101011101010";
						 when  23  =>    DADOS_AUDIO <=  "0011110101011111";
						 when  24  =>    DADOS_AUDIO <=  "0011111111001100";
						 when  25  =>    DADOS_AUDIO <=  "0100001000110010";
						 when  26  =>    DADOS_AUDIO <=  "0100010010001111";
						 when  27  =>    DADOS_AUDIO <=  "0100011011100101";
						 when  28  =>    DADOS_AUDIO <=  "0100100100110010";
						 when  29  =>    DADOS_AUDIO <=  "0100101101110110";
						 when  30  =>    DADOS_AUDIO <=  "0100110110110000";
						 when  31  =>    DADOS_AUDIO <=  "0100111111100010";
						 when  32  =>    DADOS_AUDIO <=  "0101001000001010";
						 when  33  =>    DADOS_AUDIO <=  "0101010000101000";
						 when  34  =>    DADOS_AUDIO <=  "0101011000111011";
						 when  35  =>    DADOS_AUDIO <=  "0101100001000100";
						 when  36  =>    DADOS_AUDIO <=  "0101101001000011";
						 when  37  =>    DADOS_AUDIO <=  "0101110000110111";
						 when  38  =>    DADOS_AUDIO <=  "0101111000011111";
						 when  39  =>    DADOS_AUDIO <=  "0101111111111100";
						 when  40  =>    DADOS_AUDIO <=  "0110000111001110";
						 when  41  =>    DADOS_AUDIO <=  "0110001110010011";
						 when  42  =>    DADOS_AUDIO <=  "0110010101001101";
						 when  43  =>    DADOS_AUDIO <=  "0110011011111010";
						 when  44  =>    DADOS_AUDIO <=  "0110100010011011";
						 when  45  =>    DADOS_AUDIO <=  "0110101000101111";
						 when  46  =>    DADOS_AUDIO <=  "0110101110110110";
						 when  47  =>    DADOS_AUDIO <=  "0110110100110001";
						 when  48  =>    DADOS_AUDIO <=  "0110111010011110";
						 when  49  =>    DADOS_AUDIO <=  "0110111111111110";
						 when  50  =>    DADOS_AUDIO <=  "0111000101010000";
						 when  51  =>    DADOS_AUDIO <=  "0111001010010100";
						 when  52  =>    DADOS_AUDIO <=  "0111001111001011";
						 when  53  =>    DADOS_AUDIO <=  "0111010011110011";
						 when  54  =>    DADOS_AUDIO <=  "0111011000001110";
						 when  55  =>    DADOS_AUDIO <=  "0111011100011010";
						 when  56  =>    DADOS_AUDIO <=  "0111100000011000";
						 when  57  =>    DADOS_AUDIO <=  "0111100100000111";
						 when  58  =>    DADOS_AUDIO <=  "0111100111100111";
						 when  59  =>    DADOS_AUDIO <=  "0111101010111001";
						 when  60  =>    DADOS_AUDIO <=  "0111101101111100";
						 when  61  =>    DADOS_AUDIO <=  "0111110000110000";
						 when  62  =>    DADOS_AUDIO <=  "0111110011010101";
						 when  63  =>    DADOS_AUDIO <=  "0111110101101011";
						 when  64  =>    DADOS_AUDIO <=  "0111110111110010";
						 when  65  =>    DADOS_AUDIO <=  "0111111001101001";
						 when  66  =>    DADOS_AUDIO <=  "0111111011010001";
						 when  67  =>    DADOS_AUDIO <=  "0111111100101010";
						 when  68  =>    DADOS_AUDIO <=  "0111111101110100";
						 when  69  =>    DADOS_AUDIO <=  "0111111110101110";
						 when  70  =>    DADOS_AUDIO <=  "0111111111011000";
						 when  71  =>    DADOS_AUDIO <=  "0111111111110011";
						 when  72  =>    DADOS_AUDIO <=  "0111111111111111";
						 when  73  =>    DADOS_AUDIO <=  "0111111111111011";
						 when  74  =>    DADOS_AUDIO <=  "0111111111101000";
						 when  75  =>    DADOS_AUDIO <=  "0111111111000101";
						 when  76  =>    DADOS_AUDIO <=  "0111111110010011";
						 when  77  =>    DADOS_AUDIO <=  "0111111101010001";
						 when  78  =>    DADOS_AUDIO <=  "0111111100000000";
						 when  79  =>    DADOS_AUDIO <=  "0111111010011111";
						 when  80  =>    DADOS_AUDIO <=  "0111111000101111";
						 when  81  =>    DADOS_AUDIO <=  "0111110110110000";
						 when  82  =>    DADOS_AUDIO <=  "0111110100100010";
						 when  83  =>    DADOS_AUDIO <=  "0111110010000101";
						 when  84  =>    DADOS_AUDIO <=  "0111101111011000";
						 when  85  =>    DADOS_AUDIO <=  "0111101100011101";
						 when  86  =>    DADOS_AUDIO <=  "0111101001010010";
						 when  87  =>    DADOS_AUDIO <=  "0111100101111001";
						 when  88  =>    DADOS_AUDIO <=  "0111100010010001";
						 when  89  =>    DADOS_AUDIO <=  "0111011110011011";
						 when  90  =>    DADOS_AUDIO <=  "0111011010010110";
						 when  91  =>    DADOS_AUDIO <=  "0111010110000010";
						 when  92  =>    DADOS_AUDIO <=  "0111010001100001";
						 when  93  =>    DADOS_AUDIO <=  "0111001100110001";
						 when  94  =>    DADOS_AUDIO <=  "0111000111110100";
						 when  95  =>    DADOS_AUDIO <=  "0111000010101000";
						 when  96  =>    DADOS_AUDIO <=  "0110111101001111";
						 when  97  =>    DADOS_AUDIO <=  "0110110111101001";
						 when  98  =>    DADOS_AUDIO <=  "0110110001110101";
						 when  99  =>    DADOS_AUDIO <=  "0110101011110100";
						 when  100  =>    DADOS_AUDIO <=  "0110100101100111";
						 when  101  =>    DADOS_AUDIO <=  "0110011111001100";
						 when  102  =>    DADOS_AUDIO <=  "0110011000100101";
						 when  103  =>    DADOS_AUDIO <=  "0110010001110001";
						 when  104  =>    DADOS_AUDIO <=  "0110001010110010";
						 when  105  =>    DADOS_AUDIO <=  "0110000011100110";
						 when  106  =>    DADOS_AUDIO <=  "0101111100001111";
						 when  107  =>    DADOS_AUDIO <=  "0101110100101100";
						 when  108  =>    DADOS_AUDIO <=  "0101101100111110";
						 when  109  =>    DADOS_AUDIO <=  "0101100101000101";
						 when  110  =>    DADOS_AUDIO <=  "0101011101000001";
						 when  111  =>    DADOS_AUDIO <=  "0101010100110011";
						 when  112  =>    DADOS_AUDIO <=  "0101001100011010";
						 when  113  =>    DADOS_AUDIO <=  "0101000011110111";
						 when  114  =>    DADOS_AUDIO <=  "0100111011001010";
						 when  115  =>    DADOS_AUDIO <=  "0100110010010100";
						 when  116  =>    DADOS_AUDIO <=  "0100101001010101";
						 when  117  =>    DADOS_AUDIO <=  "0100100000001100";
						 when  118  =>    DADOS_AUDIO <=  "0100010110111011";
						 when  119  =>    DADOS_AUDIO <=  "0100001101100010";
						 when  120  =>    DADOS_AUDIO <=  "0100000100000000";
						 when  121  =>    DADOS_AUDIO <=  "0011111010010110";
						 when  122  =>    DADOS_AUDIO <=  "0011110000100101";
						 when  123  =>    DADOS_AUDIO <=  "0011100110101101";
						 when  124  =>    DADOS_AUDIO <=  "0011011100101101";
						 when  125  =>    DADOS_AUDIO <=  "0011010010100111";
						 when  126  =>    DADOS_AUDIO <=  "0011001000011011";
						 when  127  =>    DADOS_AUDIO <=  "0010111110001000";
						 when  128  =>    DADOS_AUDIO <=  "0010110011110000";
						 when  129  =>    DADOS_AUDIO <=  "0010101001010010";
						 when  130  =>    DADOS_AUDIO <=  "0010011110101111";
						 when  131  =>    DADOS_AUDIO <=  "0010010100001000";
						 when  132  =>    DADOS_AUDIO <=  "0010001001011011";
						 when  133  =>    DADOS_AUDIO <=  "0001111110101011";
						 when  134  =>    DADOS_AUDIO <=  "0001110011110111";
						 when  135  =>    DADOS_AUDIO <=  "0001101000111111";
						 when  136  =>    DADOS_AUDIO <=  "0001011110000101";
						 when  137  =>    DADOS_AUDIO <=  "0001010011000111";
						 when  138  =>    DADOS_AUDIO <=  "0001001000000111";
						 when  139  =>    DADOS_AUDIO <=  "0000111101000100";
						 when  140  =>    DADOS_AUDIO <=  "0000110010000000";
						 when  141  =>    DADOS_AUDIO <=  "0000100110111011";
						 when  142  =>    DADOS_AUDIO <=  "0000011011110100";
						 when  143  =>    DADOS_AUDIO <=  "0000010000101100";
						 when  144  =>    DADOS_AUDIO <=  "0000000101100100";
						 when  145  =>    DADOS_AUDIO <=  "1111111010011100";
						 when  146  =>    DADOS_AUDIO <=  "1111101111010100";
						 when  147  =>    DADOS_AUDIO <=  "1111100100001100";
						 when  148  =>    DADOS_AUDIO <=  "1111011001000101";
						 when  149  =>    DADOS_AUDIO <=  "1111001110000000";
						 when  150  =>    DADOS_AUDIO <=  "1111000010111100";
						 when  151  =>    DADOS_AUDIO <=  "1110110111111001";
						 when  152  =>    DADOS_AUDIO <=  "1110101100111001";
						 when  153  =>    DADOS_AUDIO <=  "1110100001111011";
						 when  154  =>    DADOS_AUDIO <=  "1110010111000001";
						 when  155  =>    DADOS_AUDIO <=  "1110001100001001";
						 when  156  =>    DADOS_AUDIO <=  "1110000001010101";
						 when  157  =>    DADOS_AUDIO <=  "1101110110100101";
						 when  158  =>    DADOS_AUDIO <=  "1101101011111000";
						 when  159  =>    DADOS_AUDIO <=  "1101100001010001";
						 when  160  =>    DADOS_AUDIO <=  "1101010110101110";
						 when  161  =>    DADOS_AUDIO <=  "1101001100010000";
						 when  162  =>    DADOS_AUDIO <=  "1101000001111000";
						 when  163  =>    DADOS_AUDIO <=  "1100110111100101";
						 when  164  =>    DADOS_AUDIO <=  "1100101101011001";
						 when  165  =>    DADOS_AUDIO <=  "1100100011010011";
						 when  166  =>    DADOS_AUDIO <=  "1100011001010011";
						 when  167  =>    DADOS_AUDIO <=  "1100001111011011";
						 when  168  =>    DADOS_AUDIO <=  "1100000101101010";
						 when  169  =>    DADOS_AUDIO <=  "1011111100000000";
						 when  170  =>    DADOS_AUDIO <=  "1011110010011110";
						 when  171  =>    DADOS_AUDIO <=  "1011101001000101";
						 when  172  =>    DADOS_AUDIO <=  "1011011111110100";
						 when  173  =>    DADOS_AUDIO <=  "1011010110101011";
						 when  174  =>    DADOS_AUDIO <=  "1011001101101100";
						 when  175  =>    DADOS_AUDIO <=  "1011000100110110";
						 when  176  =>    DADOS_AUDIO <=  "1010111100001001";
						 when  177  =>    DADOS_AUDIO <=  "1010110011100110";
						 when  178  =>    DADOS_AUDIO <=  "1010101011001101";
						 when  179  =>    DADOS_AUDIO <=  "1010100010111111";
						 when  180  =>    DADOS_AUDIO <=  "1010011010111011";
						 when  181  =>    DADOS_AUDIO <=  "1010010011000010";
						 when  182  =>    DADOS_AUDIO <=  "1010001011010100";
						 when  183  =>    DADOS_AUDIO <=  "1010000011110001";
						 when  184  =>    DADOS_AUDIO <=  "1001111100011010";
						 when  185  =>    DADOS_AUDIO <=  "1001110101001110";
						 when  186  =>    DADOS_AUDIO <=  "1001101110001111";
						 when  187  =>    DADOS_AUDIO <=  "1001100111011011";
						 when  188  =>    DADOS_AUDIO <=  "1001100000110100";
						 when  189  =>    DADOS_AUDIO <=  "1001011010011001";
						 when  190  =>    DADOS_AUDIO <=  "1001010100001100";
						 when  191  =>    DADOS_AUDIO <=  "1001001110001011";
						 when  192  =>    DADOS_AUDIO <=  "1001001000010111";
						 when  193  =>    DADOS_AUDIO <=  "1001000010110001";
						 when  194  =>    DADOS_AUDIO <=  "1000111101011000";
						 when  195  =>    DADOS_AUDIO <=  "1000111000001100";
						 when  196  =>    DADOS_AUDIO <=  "1000110011001111";
						 when  197  =>    DADOS_AUDIO <=  "1000101110011111";
						 when  198  =>    DADOS_AUDIO <=  "1000101001111110";
						 when  199  =>    DADOS_AUDIO <=  "1000100101101010";
						 when  200  =>    DADOS_AUDIO <=  "1000100001100101";
						 when  201  =>    DADOS_AUDIO <=  "1000011101101111";
						 when  202  =>    DADOS_AUDIO <=  "1000011010000111";
						 when  203  =>    DADOS_AUDIO <=  "1000010110101110";
						 when  204  =>    DADOS_AUDIO <=  "1000010011100011";
						 when  205  =>    DADOS_AUDIO <=  "1000010000101000";
						 when  206  =>    DADOS_AUDIO <=  "1000001101111011";
						 when  207  =>    DADOS_AUDIO <=  "1000001011011110";
						 when  208  =>    DADOS_AUDIO <=  "1000001001010000";
						 when  209  =>    DADOS_AUDIO <=  "1000000111010001";
						 when  210  =>    DADOS_AUDIO <=  "1000000101100001";
						 when  211  =>    DADOS_AUDIO <=  "1000000100000000";
						 when  212  =>    DADOS_AUDIO <=  "1000000010101111";
						 when  213  =>    DADOS_AUDIO <=  "1000000001101101";
						 when  214  =>    DADOS_AUDIO <=  "1000000000111011";
						 when  215  =>    DADOS_AUDIO <=  "1000000000011000";
						 when  216  =>    DADOS_AUDIO <=  "1000000000000101";
						 when  217  =>    DADOS_AUDIO <=  "1000000000000001";
						 when  218  =>    DADOS_AUDIO <=  "1000000000001101";
						 when  219  =>    DADOS_AUDIO <=  "1000000000101000";
						 when  220  =>    DADOS_AUDIO <=  "1000000001010010";
						 when  221  =>    DADOS_AUDIO <=  "1000000010001100";
						 when  222  =>    DADOS_AUDIO <=  "1000000011010110";
						 when  223  =>    DADOS_AUDIO <=  "1000000100101111";
						 when  224  =>    DADOS_AUDIO <=  "1000000110010111";
						 when  225  =>    DADOS_AUDIO <=  "1000001000001110";
						 when  226  =>    DADOS_AUDIO <=  "1000001010010101";
						 when  227  =>    DADOS_AUDIO <=  "1000001100101011";
						 when  228  =>    DADOS_AUDIO <=  "1000001111010000";
						 when  229  =>    DADOS_AUDIO <=  "1000010010000100";
						 when  230  =>    DADOS_AUDIO <=  "1000010101000111";
						 when  231  =>    DADOS_AUDIO <=  "1000011000011001";
						 when  232  =>    DADOS_AUDIO <=  "1000011011111001";
						 when  233  =>    DADOS_AUDIO <=  "1000011111101000";
						 when  234  =>    DADOS_AUDIO <=  "1000100011100110";
						 when  235  =>    DADOS_AUDIO <=  "1000100111110010";
						 when  236  =>    DADOS_AUDIO <=  "1000101100001101";
						 when  237  =>    DADOS_AUDIO <=  "1000110000110101";
						 when  238  =>    DADOS_AUDIO <=  "1000110101101100";
						 when  239  =>    DADOS_AUDIO <=  "1000111010110000";
						 when  240  =>    DADOS_AUDIO <=  "1001000000000010";
						 when  241  =>    DADOS_AUDIO <=  "1001000101100010";
						 when  242  =>    DADOS_AUDIO <=  "1001001011001111";
						 when  243  =>    DADOS_AUDIO <=  "1001010001001010";
						 when  244  =>    DADOS_AUDIO <=  "1001010111010001";
						 when  245  =>    DADOS_AUDIO <=  "1001011101100101";
						 when  246  =>    DADOS_AUDIO <=  "1001100100000110";
						 when  247  =>    DADOS_AUDIO <=  "1001101010110011";
						 when  248  =>    DADOS_AUDIO <=  "1001110001101101";
						 when  249  =>    DADOS_AUDIO <=  "1001111000110010";
						 when  250  =>    DADOS_AUDIO <=  "1010000000000100";
						 when  251  =>    DADOS_AUDIO <=  "1010000111100001";
						 when  252  =>    DADOS_AUDIO <=  "1010001111001001";
						 when  253  =>    DADOS_AUDIO <=  "1010010110111101";
						 when  254  =>    DADOS_AUDIO <=  "1010011110111100";
						 when  255  =>    DADOS_AUDIO <=  "1010100111000101";
						 when  256  =>    DADOS_AUDIO <=  "1010101111011000";
						 when  257  =>    DADOS_AUDIO <=  "1010110111110110";
						 when  258  =>    DADOS_AUDIO <=  "1011000000011110";
						 when  259  =>    DADOS_AUDIO <=  "1011001001010000";
						 when  260  =>    DADOS_AUDIO <=  "1011010010001010";
						 when  261  =>    DADOS_AUDIO <=  "1011011011001110";
						 when  262  =>    DADOS_AUDIO <=  "1011100100011011";
						 when  263  =>    DADOS_AUDIO <=  "1011101101110001";
						 when  264  =>    DADOS_AUDIO <=  "1011110111001110";
						 when  265  =>    DADOS_AUDIO <=  "1100000000110100";
						 when  266  =>    DADOS_AUDIO <=  "1100001010100001";
						 when  267  =>    DADOS_AUDIO <=  "1100010100010110";
						 when  268  =>    DADOS_AUDIO <=  "1100011110010010";
						 when  269  =>    DADOS_AUDIO <=  "1100101000010101";
						 when  270  =>    DADOS_AUDIO <=  "1100110010011110";
						 when  271  =>    DADOS_AUDIO <=  "1100111100101110";
						 when  272  =>    DADOS_AUDIO <=  "1101000111000011";
						 when  273  =>    DADOS_AUDIO <=  "1101010001011110";
						 when  274  =>    DADOS_AUDIO <=  "1101011011111111";
						 when  275  =>    DADOS_AUDIO <=  "1101100110100100";
						 when  276  =>    DADOS_AUDIO <=  "1101110001001110";
						 when  277  =>    DADOS_AUDIO <=  "1101111011111100";
						 when  278  =>    DADOS_AUDIO <=  "1110000110101110";
						 when  279  =>    DADOS_AUDIO <=  "1110010001100100";
						 when  280  =>    DADOS_AUDIO <=  "1110011100011110";
						 when  281  =>    DADOS_AUDIO <=  "1110100111011010";
						 when  282  =>    DADOS_AUDIO <=  "1110110010011001";
						 when  283  =>    DADOS_AUDIO <=  "1110111101011010";
						 when  284  =>    DADOS_AUDIO <=  "1111001000011101";
						 when  285  =>    DADOS_AUDIO <=  "1111010011100010";
						 when  286  =>    DADOS_AUDIO <=  "1111011110101001";
						 when  287  =>    DADOS_AUDIO <=  "1111101001110000";
						 when  288  =>    DADOS_AUDIO <=  "1111110100111000";
						 when  289  =>    DADOS_AUDIO <=  "0000000000000000";
						 when others =>	DADOS_AUDIO <=  "0000000000000000";
					end case;
				when 6 =>
					n_pontos <= 275;
					reset <= '0';
					case aux_dados is
					    when  0  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  1  =>    DADOS_AUDIO <=  "0000001011101111";
						 when  2  =>    DADOS_AUDIO <=  "0000010111011110";
						 when  3  =>    DADOS_AUDIO <=  "0000100011001100";
						 when  4  =>    DADOS_AUDIO <=  "0000101110111001";
						 when  5  =>    DADOS_AUDIO <=  "0000111010100100";
						 when  6  =>    DADOS_AUDIO <=  "0001000110001110";
						 when  7  =>    DADOS_AUDIO <=  "0001010001110101";
						 when  8  =>    DADOS_AUDIO <=  "0001011101011001";
						 when  9  =>    DADOS_AUDIO <=  "0001101000111010";
						 when  10  =>    DADOS_AUDIO <=  "0001110100011000";
						 when  11  =>    DADOS_AUDIO <=  "0001111111110010";
						 when  12  =>    DADOS_AUDIO <=  "0010001011000111";
						 when  13  =>    DADOS_AUDIO <=  "0010010110011000";
						 when  14  =>    DADOS_AUDIO <=  "0010100001100100";
						 when  15  =>    DADOS_AUDIO <=  "0010101100101010";
						 when  16  =>    DADOS_AUDIO <=  "0010110111101010";
						 when  17  =>    DADOS_AUDIO <=  "0011000010100100";
						 when  18  =>    DADOS_AUDIO <=  "0011001101011000";
						 when  19  =>    DADOS_AUDIO <=  "0011011000000101";
						 when  20  =>    DADOS_AUDIO <=  "0011100010101010";
						 when  21  =>    DADOS_AUDIO <=  "0011101101001000";
						 when  22  =>    DADOS_AUDIO <=  "0011110111011110";
						 when  23  =>    DADOS_AUDIO <=  "0100000001101100";
						 when  24  =>    DADOS_AUDIO <=  "0100001011110001";
						 when  25  =>    DADOS_AUDIO <=  "0100010101101101";
						 when  26  =>    DADOS_AUDIO <=  "0100011111011111";
						 when  27  =>    DADOS_AUDIO <=  "0100101001001000";
						 when  28  =>    DADOS_AUDIO <=  "0100110010100111";
						 when  29  =>    DADOS_AUDIO <=  "0100111011111100";
						 when  30  =>    DADOS_AUDIO <=  "0101000101000101";
						 when  31  =>    DADOS_AUDIO <=  "0101001110000100";
						 when  32  =>    DADOS_AUDIO <=  "0101010110111000";
						 when  33  =>    DADOS_AUDIO <=  "0101011111100000";
						 when  34  =>    DADOS_AUDIO <=  "0101100111111101";
						 when  35  =>    DADOS_AUDIO <=  "0101110000001101";
						 when  36  =>    DADOS_AUDIO <=  "0101111000010001";
						 when  37  =>    DADOS_AUDIO <=  "0110000000001000";
						 when  38  =>    DADOS_AUDIO <=  "0110000111110010";
						 when  39  =>    DADOS_AUDIO <=  "0110001111001111";
						 when  40  =>    DADOS_AUDIO <=  "0110010110011111";
						 when  41  =>    DADOS_AUDIO <=  "0110011101100001";
						 when  42  =>    DADOS_AUDIO <=  "0110100100010101";
						 when  43  =>    DADOS_AUDIO <=  "0110101010111011";
						 when  44  =>    DADOS_AUDIO <=  "0110110001010011";
						 when  45  =>    DADOS_AUDIO <=  "0110110111011100";
						 when  46  =>    DADOS_AUDIO <=  "0110111101010110";
						 when  47  =>    DADOS_AUDIO <=  "0111000011000001";
						 when  48  =>    DADOS_AUDIO <=  "0111001000011101";
						 when  49  =>    DADOS_AUDIO <=  "0111001101101010";
						 when  50  =>    DADOS_AUDIO <=  "0111010010100111";
						 when  51  =>    DADOS_AUDIO <=  "0111010111010100";
						 when  52  =>    DADOS_AUDIO <=  "0111011011110010";
						 when  53  =>    DADOS_AUDIO <=  "0111011111111111";
						 when  54  =>    DADOS_AUDIO <=  "0111100011111101";
						 when  55  =>    DADOS_AUDIO <=  "0111100111101010";
						 when  56  =>    DADOS_AUDIO <=  "0111101011000111";
						 when  57  =>    DADOS_AUDIO <=  "0111101110010011";
						 when  58  =>    DADOS_AUDIO <=  "0111110001001110";
						 when  59  =>    DADOS_AUDIO <=  "0111110011111001";
						 when  60  =>    DADOS_AUDIO <=  "0111110110010011";
						 when  61  =>    DADOS_AUDIO <=  "0111111000011100";
						 when  62  =>    DADOS_AUDIO <=  "0111111010010100";
						 when  63  =>    DADOS_AUDIO <=  "0111111011111011";
						 when  64  =>    DADOS_AUDIO <=  "0111111101010001";
						 when  65  =>    DADOS_AUDIO <=  "0111111110010110";
						 when  66  =>    DADOS_AUDIO <=  "0111111111001010";
						 when  67  =>    DADOS_AUDIO <=  "0111111111101100";
						 when  68  =>    DADOS_AUDIO <=  "0111111111111101";
						 when  69  =>    DADOS_AUDIO <=  "0111111111111101";
						 when  70  =>    DADOS_AUDIO <=  "0111111111101100";
						 when  71  =>    DADOS_AUDIO <=  "0111111111001010";
						 when  72  =>    DADOS_AUDIO <=  "0111111110010110";
						 when  73  =>    DADOS_AUDIO <=  "0111111101010001";
						 when  74  =>    DADOS_AUDIO <=  "0111111011111011";
						 when  75  =>    DADOS_AUDIO <=  "0111111010010100";
						 when  76  =>    DADOS_AUDIO <=  "0111111000011100";
						 when  77  =>    DADOS_AUDIO <=  "0111110110010011";
						 when  78  =>    DADOS_AUDIO <=  "0111110011111001";
						 when  79  =>    DADOS_AUDIO <=  "0111110001001110";
						 when  80  =>    DADOS_AUDIO <=  "0111101110010011";
						 when  81  =>    DADOS_AUDIO <=  "0111101011000111";
						 when  82  =>    DADOS_AUDIO <=  "0111100111101010";
						 when  83  =>    DADOS_AUDIO <=  "0111100011111101";
						 when  84  =>    DADOS_AUDIO <=  "0111011111111111";
						 when  85  =>    DADOS_AUDIO <=  "0111011011110010";
						 when  86  =>    DADOS_AUDIO <=  "0111010111010100";
						 when  87  =>    DADOS_AUDIO <=  "0111010010100111";
						 when  88  =>    DADOS_AUDIO <=  "0111001101101010";
						 when  89  =>    DADOS_AUDIO <=  "0111001000011101";
						 when  90  =>    DADOS_AUDIO <=  "0111000011000001";
						 when  91  =>    DADOS_AUDIO <=  "0110111101010110";
						 when  92  =>    DADOS_AUDIO <=  "0110110111011100";
						 when  93  =>    DADOS_AUDIO <=  "0110110001010011";
						 when  94  =>    DADOS_AUDIO <=  "0110101010111011";
						 when  95  =>    DADOS_AUDIO <=  "0110100100010101";
						 when  96  =>    DADOS_AUDIO <=  "0110011101100001";
						 when  97  =>    DADOS_AUDIO <=  "0110010110011111";
						 when  98  =>    DADOS_AUDIO <=  "0110001111001111";
						 when  99  =>    DADOS_AUDIO <=  "0110000111110010";
						 when  100  =>    DADOS_AUDIO <=  "0110000000001000";
						 when  101  =>    DADOS_AUDIO <=  "0101111000010001";
						 when  102  =>    DADOS_AUDIO <=  "0101110000001101";
						 when  103  =>    DADOS_AUDIO <=  "0101100111111101";
						 when  104  =>    DADOS_AUDIO <=  "0101011111100000";
						 when  105  =>    DADOS_AUDIO <=  "0101010110111000";
						 when  106  =>    DADOS_AUDIO <=  "0101001110000100";
						 when  107  =>    DADOS_AUDIO <=  "0101000101000101";
						 when  108  =>    DADOS_AUDIO <=  "0100111011111100";
						 when  109  =>    DADOS_AUDIO <=  "0100110010100111";
						 when  110  =>    DADOS_AUDIO <=  "0100101001001000";
						 when  111  =>    DADOS_AUDIO <=  "0100011111011111";
						 when  112  =>    DADOS_AUDIO <=  "0100010101101101";
						 when  113  =>    DADOS_AUDIO <=  "0100001011110001";
						 when  114  =>    DADOS_AUDIO <=  "0100000001101100";
						 when  115  =>    DADOS_AUDIO <=  "0011110111011110";
						 when  116  =>    DADOS_AUDIO <=  "0011101101001000";
						 when  117  =>    DADOS_AUDIO <=  "0011100010101010";
						 when  118  =>    DADOS_AUDIO <=  "0011011000000101";
						 when  119  =>    DADOS_AUDIO <=  "0011001101011000";
						 when  120  =>    DADOS_AUDIO <=  "0011000010100100";
						 when  121  =>    DADOS_AUDIO <=  "0010110111101010";
						 when  122  =>    DADOS_AUDIO <=  "0010101100101010";
						 when  123  =>    DADOS_AUDIO <=  "0010100001100100";
						 when  124  =>    DADOS_AUDIO <=  "0010010110011000";
						 when  125  =>    DADOS_AUDIO <=  "0010001011000111";
						 when  126  =>    DADOS_AUDIO <=  "0001111111110010";
						 when  127  =>    DADOS_AUDIO <=  "0001110100011000";
						 when  128  =>    DADOS_AUDIO <=  "0001101000111010";
						 when  129  =>    DADOS_AUDIO <=  "0001011101011001";
						 when  130  =>    DADOS_AUDIO <=  "0001010001110101";
						 when  131  =>    DADOS_AUDIO <=  "0001000110001110";
						 when  132  =>    DADOS_AUDIO <=  "0000111010100100";
						 when  133  =>    DADOS_AUDIO <=  "0000101110111001";
						 when  134  =>    DADOS_AUDIO <=  "0000100011001100";
						 when  135  =>    DADOS_AUDIO <=  "0000010111011110";
						 when  136  =>    DADOS_AUDIO <=  "0000001011101111";
						 when  137  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  138  =>    DADOS_AUDIO <=  "1111110100010001";
						 when  139  =>    DADOS_AUDIO <=  "1111101000100010";
						 when  140  =>    DADOS_AUDIO <=  "1111011100110100";
						 when  141  =>    DADOS_AUDIO <=  "1111010001000111";
						 when  142  =>    DADOS_AUDIO <=  "1111000101011100";
						 when  143  =>    DADOS_AUDIO <=  "1110111001110010";
						 when  144  =>    DADOS_AUDIO <=  "1110101110001011";
						 when  145  =>    DADOS_AUDIO <=  "1110100010100111";
						 when  146  =>    DADOS_AUDIO <=  "1110010111000110";
						 when  147  =>    DADOS_AUDIO <=  "1110001011101000";
						 when  148  =>    DADOS_AUDIO <=  "1110000000001110";
						 when  149  =>    DADOS_AUDIO <=  "1101110100111001";
						 when  150  =>    DADOS_AUDIO <=  "1101101001101000";
						 when  151  =>    DADOS_AUDIO <=  "1101011110011100";
						 when  152  =>    DADOS_AUDIO <=  "1101010011010110";
						 when  153  =>    DADOS_AUDIO <=  "1101001000010110";
						 when  154  =>    DADOS_AUDIO <=  "1100111101011100";
						 when  155  =>    DADOS_AUDIO <=  "1100110010101000";
						 when  156  =>    DADOS_AUDIO <=  "1100100111111011";
						 when  157  =>    DADOS_AUDIO <=  "1100011101010110";
						 when  158  =>    DADOS_AUDIO <=  "1100010010111000";
						 when  159  =>    DADOS_AUDIO <=  "1100001000100010";
						 when  160  =>    DADOS_AUDIO <=  "1011111110010100";
						 when  161  =>    DADOS_AUDIO <=  "1011110100001111";
						 when  162  =>    DADOS_AUDIO <=  "1011101010010011";
						 when  163  =>    DADOS_AUDIO <=  "1011100000100001";
						 when  164  =>    DADOS_AUDIO <=  "1011010110111000";
						 when  165  =>    DADOS_AUDIO <=  "1011001101011001";
						 when  166  =>    DADOS_AUDIO <=  "1011000100000100";
						 when  167  =>    DADOS_AUDIO <=  "1010111010111011";
						 when  168  =>    DADOS_AUDIO <=  "1010110001111100";
						 when  169  =>    DADOS_AUDIO <=  "1010101001001000";
						 when  170  =>    DADOS_AUDIO <=  "1010100000100000";
						 when  171  =>    DADOS_AUDIO <=  "1010011000000011";
						 when  172  =>    DADOS_AUDIO <=  "1010001111110011";
						 when  173  =>    DADOS_AUDIO <=  "1010000111101111";
						 when  174  =>    DADOS_AUDIO <=  "1001111111111000";
						 when  175  =>    DADOS_AUDIO <=  "1001111000001110";
						 when  176  =>    DADOS_AUDIO <=  "1001110000110001";
						 when  177  =>    DADOS_AUDIO <=  "1001101001100001";
						 when  178  =>    DADOS_AUDIO <=  "1001100010011111";
						 when  179  =>    DADOS_AUDIO <=  "1001011011101011";
						 when  180  =>    DADOS_AUDIO <=  "1001010101000101";
						 when  181  =>    DADOS_AUDIO <=  "1001001110101101";
						 when  182  =>    DADOS_AUDIO <=  "1001001000100100";
						 when  183  =>    DADOS_AUDIO <=  "1001000010101010";
						 when  184  =>    DADOS_AUDIO <=  "1000111100111111";
						 when  185  =>    DADOS_AUDIO <=  "1000110111100011";
						 when  186  =>    DADOS_AUDIO <=  "1000110010010110";
						 when  187  =>    DADOS_AUDIO <=  "1000101101011001";
						 when  188  =>    DADOS_AUDIO <=  "1000101000101100";
						 when  189  =>    DADOS_AUDIO <=  "1000100100001110";
						 when  190  =>    DADOS_AUDIO <=  "1000100000000001";
						 when  191  =>    DADOS_AUDIO <=  "1000011100000011";
						 when  192  =>    DADOS_AUDIO <=  "1000011000010110";
						 when  193  =>    DADOS_AUDIO <=  "1000010100111001";
						 when  194  =>    DADOS_AUDIO <=  "1000010001101101";
						 when  195  =>    DADOS_AUDIO <=  "1000001110110010";
						 when  196  =>    DADOS_AUDIO <=  "1000001100000111";
						 when  197  =>    DADOS_AUDIO <=  "1000001001101101";
						 when  198  =>    DADOS_AUDIO <=  "1000000111100100";
						 when  199  =>    DADOS_AUDIO <=  "1000000101101100";
						 when  200  =>    DADOS_AUDIO <=  "1000000100000101";
						 when  201  =>    DADOS_AUDIO <=  "1000000010101111";
						 when  202  =>    DADOS_AUDIO <=  "1000000001101010";
						 when  203  =>    DADOS_AUDIO <=  "1000000000110110";
						 when  204  =>    DADOS_AUDIO <=  "1000000000010100";
						 when  205  =>    DADOS_AUDIO <=  "1000000000000011";
						 when  206  =>    DADOS_AUDIO <=  "1000000000000011";
						 when  207  =>    DADOS_AUDIO <=  "1000000000010100";
						 when  208  =>    DADOS_AUDIO <=  "1000000000110110";
						 when  209  =>    DADOS_AUDIO <=  "1000000001101010";
						 when  210  =>    DADOS_AUDIO <=  "1000000010101111";
						 when  211  =>    DADOS_AUDIO <=  "1000000100000101";
						 when  212  =>    DADOS_AUDIO <=  "1000000101101100";
						 when  213  =>    DADOS_AUDIO <=  "1000000111100100";
						 when  214  =>    DADOS_AUDIO <=  "1000001001101101";
						 when  215  =>    DADOS_AUDIO <=  "1000001100000111";
						 when  216  =>    DADOS_AUDIO <=  "1000001110110010";
						 when  217  =>    DADOS_AUDIO <=  "1000010001101101";
						 when  218  =>    DADOS_AUDIO <=  "1000010100111001";
						 when  219  =>    DADOS_AUDIO <=  "1000011000010110";
						 when  220  =>    DADOS_AUDIO <=  "1000011100000011";
						 when  221  =>    DADOS_AUDIO <=  "1000100000000001";
						 when  222  =>    DADOS_AUDIO <=  "1000100100001110";
						 when  223  =>    DADOS_AUDIO <=  "1000101000101100";
						 when  224  =>    DADOS_AUDIO <=  "1000101101011001";
						 when  225  =>    DADOS_AUDIO <=  "1000110010010110";
						 when  226  =>    DADOS_AUDIO <=  "1000110111100011";
						 when  227  =>    DADOS_AUDIO <=  "1000111100111111";
						 when  228  =>    DADOS_AUDIO <=  "1001000010101010";
						 when  229  =>    DADOS_AUDIO <=  "1001001000100100";
						 when  230  =>    DADOS_AUDIO <=  "1001001110101101";
						 when  231  =>    DADOS_AUDIO <=  "1001010101000101";
						 when  232  =>    DADOS_AUDIO <=  "1001011011101011";
						 when  233  =>    DADOS_AUDIO <=  "1001100010011111";
						 when  234  =>    DADOS_AUDIO <=  "1001101001100001";
						 when  235  =>    DADOS_AUDIO <=  "1001110000110001";
						 when  236  =>    DADOS_AUDIO <=  "1001111000001110";
						 when  237  =>    DADOS_AUDIO <=  "1001111111111000";
						 when  238  =>    DADOS_AUDIO <=  "1010000111101111";
						 when  239  =>    DADOS_AUDIO <=  "1010001111110011";
						 when  240  =>    DADOS_AUDIO <=  "1010011000000011";
						 when  241  =>    DADOS_AUDIO <=  "1010100000100000";
						 when  242  =>    DADOS_AUDIO <=  "1010101001001000";
						 when  243  =>    DADOS_AUDIO <=  "1010110001111100";
						 when  244  =>    DADOS_AUDIO <=  "1010111010111011";
						 when  245  =>    DADOS_AUDIO <=  "1011000100000100";
						 when  246  =>    DADOS_AUDIO <=  "1011001101011001";
						 when  247  =>    DADOS_AUDIO <=  "1011010110111000";
						 when  248  =>    DADOS_AUDIO <=  "1011100000100001";
						 when  249  =>    DADOS_AUDIO <=  "1011101010010011";
						 when  250  =>    DADOS_AUDIO <=  "1011110100001111";
						 when  251  =>    DADOS_AUDIO <=  "1011111110010100";
						 when  252  =>    DADOS_AUDIO <=  "1100001000100010";
						 when  253  =>    DADOS_AUDIO <=  "1100010010111000";
						 when  254  =>    DADOS_AUDIO <=  "1100011101010110";
						 when  255  =>    DADOS_AUDIO <=  "1100100111111011";
						 when  256  =>    DADOS_AUDIO <=  "1100110010101000";
						 when  257  =>    DADOS_AUDIO <=  "1100111101011100";
						 when  258  =>    DADOS_AUDIO <=  "1101001000010110";
						 when  259  =>    DADOS_AUDIO <=  "1101010011010110";
						 when  260  =>    DADOS_AUDIO <=  "1101011110011100";
						 when  261  =>    DADOS_AUDIO <=  "1101101001101000";
						 when  262  =>    DADOS_AUDIO <=  "1101110100111001";
						 when  263  =>    DADOS_AUDIO <=  "1110000000001110";
						 when  264  =>    DADOS_AUDIO <=  "1110001011101000";
						 when  265  =>    DADOS_AUDIO <=  "1110010111000110";
						 when  266  =>    DADOS_AUDIO <=  "1110100010100111";
						 when  267  =>    DADOS_AUDIO <=  "1110101110001011";
						 when  268  =>    DADOS_AUDIO <=  "1110111001110010";
						 when  269  =>    DADOS_AUDIO <=  "1111000101011100";
						 when  270  =>    DADOS_AUDIO <=  "1111010001000111";
						 when  271  =>    DADOS_AUDIO <=  "1111011100110100";
						 when  272  =>    DADOS_AUDIO <=  "1111101000100010";
						 when  273  =>    DADOS_AUDIO <=  "1111110100010001";
						 when  274  =>    DADOS_AUDIO <=  "0000000000000000";
						 when others =>	DADOS_AUDIO <=  "0000000000000000";
					end case;
				when 7 =>
					n_pontos <= 259;
					reset <= '0';
					case aux_dados is
					    when  0  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  1  =>    DADOS_AUDIO <=  "0000001100011101";
						 when  2  =>    DADOS_AUDIO <=  "0000011000111011";
						 when  3  =>    DADOS_AUDIO <=  "0000100101010111";
						 when  4  =>    DADOS_AUDIO <=  "0000110001110011";
						 when  5  =>    DADOS_AUDIO <=  "0000111110001100";
						 when  6  =>    DADOS_AUDIO <=  "0001001010100011";
						 when  7  =>    DADOS_AUDIO <=  "0001010110110111";
						 when  8  =>    DADOS_AUDIO <=  "0001100011000111";
						 when  9  =>    DADOS_AUDIO <=  "0001101111010100";
						 when  10  =>    DADOS_AUDIO <=  "0001111011011101";
						 when  11  =>    DADOS_AUDIO <=  "0010000111100001";
						 when  12  =>    DADOS_AUDIO <=  "0010010011100000";
						 when  13  =>    DADOS_AUDIO <=  "0010011111011001";
						 when  14  =>    DADOS_AUDIO <=  "0010101011001100";
						 when  15  =>    DADOS_AUDIO <=  "0010110110111001";
						 when  16  =>    DADOS_AUDIO <=  "0011000010011111";
						 when  17  =>    DADOS_AUDIO <=  "0011001101111101";
						 when  18  =>    DADOS_AUDIO <=  "0011011001010100";
						 when  19  =>    DADOS_AUDIO <=  "0011100100100010";
						 when  20  =>    DADOS_AUDIO <=  "0011101111101000";
						 when  21  =>    DADOS_AUDIO <=  "0011111010100101";
						 when  22  =>    DADOS_AUDIO <=  "0100000101011000";
						 when  23  =>    DADOS_AUDIO <=  "0100010000000001";
						 when  24  =>    DADOS_AUDIO <=  "0100011010100000";
						 when  25  =>    DADOS_AUDIO <=  "0100100100110100";
						 when  26  =>    DADOS_AUDIO <=  "0100101110111101";
						 when  27  =>    DADOS_AUDIO <=  "0100111000111010";
						 when  28  =>    DADOS_AUDIO <=  "0101000010101100";
						 when  29  =>    DADOS_AUDIO <=  "0101001100010001";
						 when  30  =>    DADOS_AUDIO <=  "0101010101101010";
						 when  31  =>    DADOS_AUDIO <=  "0101011110110110";
						 when  32  =>    DADOS_AUDIO <=  "0101100111110100";
						 when  33  =>    DADOS_AUDIO <=  "0101110000100101";
						 when  34  =>    DADOS_AUDIO <=  "0101111001001000";
						 when  35  =>    DADOS_AUDIO <=  "0110000001011101";
						 when  36  =>    DADOS_AUDIO <=  "0110001001100011";
						 when  37  =>    DADOS_AUDIO <=  "0110010001011001";
						 when  38  =>    DADOS_AUDIO <=  "0110011001000001";
						 when  39  =>    DADOS_AUDIO <=  "0110100000011001";
						 when  40  =>    DADOS_AUDIO <=  "0110100111100010";
						 when  41  =>    DADOS_AUDIO <=  "0110101110011010";
						 when  42  =>    DADOS_AUDIO <=  "0110110101000010";
						 when  43  =>    DADOS_AUDIO <=  "0110111011011001";
						 when  44  =>    DADOS_AUDIO <=  "0111000001100000";
						 when  45  =>    DADOS_AUDIO <=  "0111000111010101";
						 when  46  =>    DADOS_AUDIO <=  "0111001100111010";
						 when  47  =>    DADOS_AUDIO <=  "0111010010001100";
						 when  48  =>    DADOS_AUDIO <=  "0111010111001101";
						 when  49  =>    DADOS_AUDIO <=  "0111011011111101";
						 when  50  =>    DADOS_AUDIO <=  "0111100000011010";
						 when  51  =>    DADOS_AUDIO <=  "0111100100100100";
						 when  52  =>    DADOS_AUDIO <=  "0111101000011101";
						 when  53  =>    DADOS_AUDIO <=  "0111101100000011";
						 when  54  =>    DADOS_AUDIO <=  "0111101111010110";
						 when  55  =>    DADOS_AUDIO <=  "0111110010010110";
						 when  56  =>    DADOS_AUDIO <=  "0111110101000100";
						 when  57  =>    DADOS_AUDIO <=  "0111110111011110";
						 when  58  =>    DADOS_AUDIO <=  "0111111001100110";
						 when  59  =>    DADOS_AUDIO <=  "0111111011011010";
						 when  60  =>    DADOS_AUDIO <=  "0111111100111011";
						 when  61  =>    DADOS_AUDIO <=  "0111111110001001";
						 when  62  =>    DADOS_AUDIO <=  "0111111111000011";
						 when  63  =>    DADOS_AUDIO <=  "0111111111101010";
						 when  64  =>    DADOS_AUDIO <=  "0111111111111101";
						 when  65  =>    DADOS_AUDIO <=  "0111111111111101";
						 when  66  =>    DADOS_AUDIO <=  "0111111111101010";
						 when  67  =>    DADOS_AUDIO <=  "0111111111000011";
						 when  68  =>    DADOS_AUDIO <=  "0111111110001001";
						 when  69  =>    DADOS_AUDIO <=  "0111111100111011";
						 when  70  =>    DADOS_AUDIO <=  "0111111011011010";
						 when  71  =>    DADOS_AUDIO <=  "0111111001100110";
						 when  72  =>    DADOS_AUDIO <=  "0111110111011110";
						 when  73  =>    DADOS_AUDIO <=  "0111110101000100";
						 when  74  =>    DADOS_AUDIO <=  "0111110010010110";
						 when  75  =>    DADOS_AUDIO <=  "0111101111010110";
						 when  76  =>    DADOS_AUDIO <=  "0111101100000011";
						 when  77  =>    DADOS_AUDIO <=  "0111101000011101";
						 when  78  =>    DADOS_AUDIO <=  "0111100100100100";
						 when  79  =>    DADOS_AUDIO <=  "0111100000011010";
						 when  80  =>    DADOS_AUDIO <=  "0111011011111101";
						 when  81  =>    DADOS_AUDIO <=  "0111010111001101";
						 when  82  =>    DADOS_AUDIO <=  "0111010010001100";
						 when  83  =>    DADOS_AUDIO <=  "0111001100111010";
						 when  84  =>    DADOS_AUDIO <=  "0111000111010101";
						 when  85  =>    DADOS_AUDIO <=  "0111000001100000";
						 when  86  =>    DADOS_AUDIO <=  "0110111011011001";
						 when  87  =>    DADOS_AUDIO <=  "0110110101000010";
						 when  88  =>    DADOS_AUDIO <=  "0110101110011010";
						 when  89  =>    DADOS_AUDIO <=  "0110100111100010";
						 when  90  =>    DADOS_AUDIO <=  "0110100000011001";
						 when  91  =>    DADOS_AUDIO <=  "0110011001000001";
						 when  92  =>    DADOS_AUDIO <=  "0110010001011001";
						 when  93  =>    DADOS_AUDIO <=  "0110001001100011";
						 when  94  =>    DADOS_AUDIO <=  "0110000001011101";
						 when  95  =>    DADOS_AUDIO <=  "0101111001001000";
						 when  96  =>    DADOS_AUDIO <=  "0101110000100101";
						 when  97  =>    DADOS_AUDIO <=  "0101100111110100";
						 when  98  =>    DADOS_AUDIO <=  "0101011110110110";
						 when  99  =>    DADOS_AUDIO <=  "0101010101101010";
						 when  100  =>    DADOS_AUDIO <=  "0101001100010001";
						 when  101  =>    DADOS_AUDIO <=  "0101000010101100";
						 when  102  =>    DADOS_AUDIO <=  "0100111000111010";
						 when  103  =>    DADOS_AUDIO <=  "0100101110111101";
						 when  104  =>    DADOS_AUDIO <=  "0100100100110100";
						 when  105  =>    DADOS_AUDIO <=  "0100011010100000";
						 when  106  =>    DADOS_AUDIO <=  "0100010000000001";
						 when  107  =>    DADOS_AUDIO <=  "0100000101011000";
						 when  108  =>    DADOS_AUDIO <=  "0011111010100101";
						 when  109  =>    DADOS_AUDIO <=  "0011101111101000";
						 when  110  =>    DADOS_AUDIO <=  "0011100100100010";
						 when  111  =>    DADOS_AUDIO <=  "0011011001010100";
						 when  112  =>    DADOS_AUDIO <=  "0011001101111101";
						 when  113  =>    DADOS_AUDIO <=  "0011000010011111";
						 when  114  =>    DADOS_AUDIO <=  "0010110110111001";
						 when  115  =>    DADOS_AUDIO <=  "0010101011001100";
						 when  116  =>    DADOS_AUDIO <=  "0010011111011001";
						 when  117  =>    DADOS_AUDIO <=  "0010010011100000";
						 when  118  =>    DADOS_AUDIO <=  "0010000111100001";
						 when  119  =>    DADOS_AUDIO <=  "0001111011011101";
						 when  120  =>    DADOS_AUDIO <=  "0001101111010100";
						 when  121  =>    DADOS_AUDIO <=  "0001100011000111";
						 when  122  =>    DADOS_AUDIO <=  "0001010110110111";
						 when  123  =>    DADOS_AUDIO <=  "0001001010100011";
						 when  124  =>    DADOS_AUDIO <=  "0000111110001100";
						 when  125  =>    DADOS_AUDIO <=  "0000110001110011";
						 when  126  =>    DADOS_AUDIO <=  "0000100101010111";
						 when  127  =>    DADOS_AUDIO <=  "0000011000111011";
						 when  128  =>    DADOS_AUDIO <=  "0000001100011101";
						 when  129  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  130  =>    DADOS_AUDIO <=  "1111110011100011";
						 when  131  =>    DADOS_AUDIO <=  "1111100111000101";
						 when  132  =>    DADOS_AUDIO <=  "1111011010101001";
						 when  133  =>    DADOS_AUDIO <=  "1111001110001101";
						 when  134  =>    DADOS_AUDIO <=  "1111000001110100";
						 when  135  =>    DADOS_AUDIO <=  "1110110101011101";
						 when  136  =>    DADOS_AUDIO <=  "1110101001001001";
						 when  137  =>    DADOS_AUDIO <=  "1110011100111001";
						 when  138  =>    DADOS_AUDIO <=  "1110010000101100";
						 when  139  =>    DADOS_AUDIO <=  "1110000100100011";
						 when  140  =>    DADOS_AUDIO <=  "1101111000011111";
						 when  141  =>    DADOS_AUDIO <=  "1101101100100000";
						 when  142  =>    DADOS_AUDIO <=  "1101100000100111";
						 when  143  =>    DADOS_AUDIO <=  "1101010100110100";
						 when  144  =>    DADOS_AUDIO <=  "1101001001000111";
						 when  145  =>    DADOS_AUDIO <=  "1100111101100001";
						 when  146  =>    DADOS_AUDIO <=  "1100110010000011";
						 when  147  =>    DADOS_AUDIO <=  "1100100110101100";
						 when  148  =>    DADOS_AUDIO <=  "1100011011011110";
						 when  149  =>    DADOS_AUDIO <=  "1100010000011000";
						 when  150  =>    DADOS_AUDIO <=  "1100000101011011";
						 when  151  =>    DADOS_AUDIO <=  "1011111010101000";
						 when  152  =>    DADOS_AUDIO <=  "1011101111111111";
						 when  153  =>    DADOS_AUDIO <=  "1011100101100000";
						 when  154  =>    DADOS_AUDIO <=  "1011011011001100";
						 when  155  =>    DADOS_AUDIO <=  "1011010001000011";
						 when  156  =>    DADOS_AUDIO <=  "1011000111000110";
						 when  157  =>    DADOS_AUDIO <=  "1010111101010100";
						 when  158  =>    DADOS_AUDIO <=  "1010110011101111";
						 when  159  =>    DADOS_AUDIO <=  "1010101010010110";
						 when  160  =>    DADOS_AUDIO <=  "1010100001001010";
						 when  161  =>    DADOS_AUDIO <=  "1010011000001100";
						 when  162  =>    DADOS_AUDIO <=  "1010001111011011";
						 when  163  =>    DADOS_AUDIO <=  "1010000110111000";
						 when  164  =>    DADOS_AUDIO <=  "1001111110100011";
						 when  165  =>    DADOS_AUDIO <=  "1001110110011101";
						 when  166  =>    DADOS_AUDIO <=  "1001101110100111";
						 when  167  =>    DADOS_AUDIO <=  "1001100110111111";
						 when  168  =>    DADOS_AUDIO <=  "1001011111100111";
						 when  169  =>    DADOS_AUDIO <=  "1001011000011110";
						 when  170  =>    DADOS_AUDIO <=  "1001010001100110";
						 when  171  =>    DADOS_AUDIO <=  "1001001010111110";
						 when  172  =>    DADOS_AUDIO <=  "1001000100100111";
						 when  173  =>    DADOS_AUDIO <=  "1000111110100000";
						 when  174  =>    DADOS_AUDIO <=  "1000111000101011";
						 when  175  =>    DADOS_AUDIO <=  "1000110011000110";
						 when  176  =>    DADOS_AUDIO <=  "1000101101110100";
						 when  177  =>    DADOS_AUDIO <=  "1000101000110011";
						 when  178  =>    DADOS_AUDIO <=  "1000100100000011";
						 when  179  =>    DADOS_AUDIO <=  "1000011111100110";
						 when  180  =>    DADOS_AUDIO <=  "1000011011011100";
						 when  181  =>    DADOS_AUDIO <=  "1000010111100011";
						 when  182  =>    DADOS_AUDIO <=  "1000010011111101";
						 when  183  =>    DADOS_AUDIO <=  "1000010000101010";
						 when  184  =>    DADOS_AUDIO <=  "1000001101101010";
						 when  185  =>    DADOS_AUDIO <=  "1000001010111100";
						 when  186  =>    DADOS_AUDIO <=  "1000001000100010";
						 when  187  =>    DADOS_AUDIO <=  "1000000110011010";
						 when  188  =>    DADOS_AUDIO <=  "1000000100100110";
						 when  189  =>    DADOS_AUDIO <=  "1000000011000101";
						 when  190  =>    DADOS_AUDIO <=  "1000000001110111";
						 when  191  =>    DADOS_AUDIO <=  "1000000000111101";
						 when  192  =>    DADOS_AUDIO <=  "1000000000010110";
						 when  193  =>    DADOS_AUDIO <=  "1000000000000011";
						 when  194  =>    DADOS_AUDIO <=  "1000000000000011";
						 when  195  =>    DADOS_AUDIO <=  "1000000000010110";
						 when  196  =>    DADOS_AUDIO <=  "1000000000111101";
						 when  197  =>    DADOS_AUDIO <=  "1000000001110111";
						 when  198  =>    DADOS_AUDIO <=  "1000000011000101";
						 when  199  =>    DADOS_AUDIO <=  "1000000100100110";
						 when  200  =>    DADOS_AUDIO <=  "1000000110011010";
						 when  201  =>    DADOS_AUDIO <=  "1000001000100010";
						 when  202  =>    DADOS_AUDIO <=  "1000001010111100";
						 when  203  =>    DADOS_AUDIO <=  "1000001101101010";
						 when  204  =>    DADOS_AUDIO <=  "1000010000101010";
						 when  205  =>    DADOS_AUDIO <=  "1000010011111101";
						 when  206  =>    DADOS_AUDIO <=  "1000010111100011";
						 when  207  =>    DADOS_AUDIO <=  "1000011011011100";
						 when  208  =>    DADOS_AUDIO <=  "1000011111100110";
						 when  209  =>    DADOS_AUDIO <=  "1000100100000011";
						 when  210  =>    DADOS_AUDIO <=  "1000101000110011";
						 when  211  =>    DADOS_AUDIO <=  "1000101101110100";
						 when  212  =>    DADOS_AUDIO <=  "1000110011000110";
						 when  213  =>    DADOS_AUDIO <=  "1000111000101011";
						 when  214  =>    DADOS_AUDIO <=  "1000111110100000";
						 when  215  =>    DADOS_AUDIO <=  "1001000100100111";
						 when  216  =>    DADOS_AUDIO <=  "1001001010111110";
						 when  217  =>    DADOS_AUDIO <=  "1001010001100110";
						 when  218  =>    DADOS_AUDIO <=  "1001011000011110";
						 when  219  =>    DADOS_AUDIO <=  "1001011111100111";
						 when  220  =>    DADOS_AUDIO <=  "1001100110111111";
						 when  221  =>    DADOS_AUDIO <=  "1001101110100111";
						 when  222  =>    DADOS_AUDIO <=  "1001110110011101";
						 when  223  =>    DADOS_AUDIO <=  "1001111110100011";
						 when  224  =>    DADOS_AUDIO <=  "1010000110111000";
						 when  225  =>    DADOS_AUDIO <=  "1010001111011011";
						 when  226  =>    DADOS_AUDIO <=  "1010011000001100";
						 when  227  =>    DADOS_AUDIO <=  "1010100001001010";
						 when  228  =>    DADOS_AUDIO <=  "1010101010010110";
						 when  229  =>    DADOS_AUDIO <=  "1010110011101111";
						 when  230  =>    DADOS_AUDIO <=  "1010111101010100";
						 when  231  =>    DADOS_AUDIO <=  "1011000111000110";
						 when  232  =>    DADOS_AUDIO <=  "1011010001000011";
						 when  233  =>    DADOS_AUDIO <=  "1011011011001100";
						 when  234  =>    DADOS_AUDIO <=  "1011100101100000";
						 when  235  =>    DADOS_AUDIO <=  "1011101111111111";
						 when  236  =>    DADOS_AUDIO <=  "1011111010101000";
						 when  237  =>    DADOS_AUDIO <=  "1100000101011011";
						 when  238  =>    DADOS_AUDIO <=  "1100010000011000";
						 when  239  =>    DADOS_AUDIO <=  "1100011011011110";
						 when  240  =>    DADOS_AUDIO <=  "1100100110101100";
						 when  241  =>    DADOS_AUDIO <=  "1100110010000011";
						 when  242  =>    DADOS_AUDIO <=  "1100111101100001";
						 when  243  =>    DADOS_AUDIO <=  "1101001001000111";
						 when  244  =>    DADOS_AUDIO <=  "1101010100110100";
						 when  245  =>    DADOS_AUDIO <=  "1101100000100111";
						 when  246  =>    DADOS_AUDIO <=  "1101101100100000";
						 when  247  =>    DADOS_AUDIO <=  "1101111000011111";
						 when  248  =>    DADOS_AUDIO <=  "1110000100100011";
						 when  249  =>    DADOS_AUDIO <=  "1110010000101100";
						 when  250  =>    DADOS_AUDIO <=  "1110011100111001";
						 when  251  =>    DADOS_AUDIO <=  "1110101001001001";
						 when  252  =>    DADOS_AUDIO <=  "1110110101011101";
						 when  253  =>    DADOS_AUDIO <=  "1111000001110100";
						 when  254  =>    DADOS_AUDIO <=  "1111001110001101";
						 when  255  =>    DADOS_AUDIO <=  "1111011010101001";
						 when  256  =>    DADOS_AUDIO <=  "1111100111000101";
						 when  257  =>    DADOS_AUDIO <=  "1111110011100011";
						 when  258  =>    DADOS_AUDIO <=  "0000000000000000";
						 when others =>	DADOS_AUDIO <=  "0000000000000000";
					end case;
				when 8 =>
					n_pontos <= 244;
					reset <= '0';
					case aux_dados is
					    when  0  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  1  =>    DADOS_AUDIO <=  "0000001101001111";
						 when  2  =>    DADOS_AUDIO <=  "0000011010011101";
						 when  3  =>    DADOS_AUDIO <=  "0000100111101011";
						 when  4  =>    DADOS_AUDIO <=  "0000110100110111";
						 when  5  =>    DADOS_AUDIO <=  "0001000010000000";
						 when  6  =>    DADOS_AUDIO <=  "0001001111000111";
						 when  7  =>    DADOS_AUDIO <=  "0001011100001010";
						 when  8  =>    DADOS_AUDIO <=  "0001101001001001";
						 when  9  =>    DADOS_AUDIO <=  "0001110110000100";
						 when  10  =>    DADOS_AUDIO <=  "0010000010111010";
						 when  11  =>    DADOS_AUDIO <=  "0010001111101010";
						 when  12  =>    DADOS_AUDIO <=  "0010011100010100";
						 when  13  =>    DADOS_AUDIO <=  "0010101000111000";
						 when  14  =>    DADOS_AUDIO <=  "0010110101010100";
						 when  15  =>    DADOS_AUDIO <=  "0011000001101000";
						 when  16  =>    DADOS_AUDIO <=  "0011001101110100";
						 when  17  =>    DADOS_AUDIO <=  "0011011001111000";
						 when  18  =>    DADOS_AUDIO <=  "0011100101110010";
						 when  19  =>    DADOS_AUDIO <=  "0011110001100010";
						 when  20  =>    DADOS_AUDIO <=  "0011111101001000";
						 when  21  =>    DADOS_AUDIO <=  "0100001000100011";
						 when  22  =>    DADOS_AUDIO <=  "0100010011110010";
						 when  23  =>    DADOS_AUDIO <=  "0100011110110110";
						 when  24  =>    DADOS_AUDIO <=  "0100101001101110";
						 when  25  =>    DADOS_AUDIO <=  "0100110100011001";
						 when  26  =>    DADOS_AUDIO <=  "0100111110110110";
						 when  27  =>    DADOS_AUDIO <=  "0101001001000110";
						 when  28  =>    DADOS_AUDIO <=  "0101010011001000";
						 when  29  =>    DADOS_AUDIO <=  "0101011100111100";
						 when  30  =>    DADOS_AUDIO <=  "0101100110100000";
						 when  31  =>    DADOS_AUDIO <=  "0101101111110101";
						 when  32  =>    DADOS_AUDIO <=  "0101111000111011";
						 when  33  =>    DADOS_AUDIO <=  "0110000001110000";
						 when  34  =>    DADOS_AUDIO <=  "0110001010010101";
						 when  35  =>    DADOS_AUDIO <=  "0110010010101001";
						 when  36  =>    DADOS_AUDIO <=  "0110011010101011";
						 when  37  =>    DADOS_AUDIO <=  "0110100010011101";
						 when  38  =>    DADOS_AUDIO <=  "0110101001111100";
						 when  39  =>    DADOS_AUDIO <=  "0110110001001001";
						 when  40  =>    DADOS_AUDIO <=  "0110111000000011";
						 when  41  =>    DADOS_AUDIO <=  "0110111110101011";
						 when  42  =>    DADOS_AUDIO <=  "0111000100111111";
						 when  43  =>    DADOS_AUDIO <=  "0111001011000001";
						 when  44  =>    DADOS_AUDIO <=  "0111010000101110";
						 when  45  =>    DADOS_AUDIO <=  "0111010110001000";
						 when  46  =>    DADOS_AUDIO <=  "0111011011001101";
						 when  47  =>    DADOS_AUDIO <=  "0111011111111110";
						 when  48  =>    DADOS_AUDIO <=  "0111100100011011";
						 when  49  =>    DADOS_AUDIO <=  "0111101000100011";
						 when  50  =>    DADOS_AUDIO <=  "0111101100010110";
						 when  51  =>    DADOS_AUDIO <=  "0111101111110100";
						 when  52  =>    DADOS_AUDIO <=  "0111110010111100";
						 when  53  =>    DADOS_AUDIO <=  "0111110101110000";
						 when  54  =>    DADOS_AUDIO <=  "0111111000001110";
						 when  55  =>    DADOS_AUDIO <=  "0111111010010110";
						 when  56  =>    DADOS_AUDIO <=  "0111111100001001";
						 when  57  =>    DADOS_AUDIO <=  "0111111101100110";
						 when  58  =>    DADOS_AUDIO <=  "0111111110101101";
						 when  59  =>    DADOS_AUDIO <=  "0111111111011110";
						 when  60  =>    DADOS_AUDIO <=  "0111111111111001";
						 when  61  =>    DADOS_AUDIO <=  "0111111111111111";
						 when  62  =>    DADOS_AUDIO <=  "0111111111101110";
						 when  63  =>    DADOS_AUDIO <=  "0111111111001000";
						 when  64  =>    DADOS_AUDIO <=  "0111111110001100";
						 when  65  =>    DADOS_AUDIO <=  "0111111100111010";
						 when  66  =>    DADOS_AUDIO <=  "0111111011010010";
						 when  67  =>    DADOS_AUDIO <=  "0111111001010101";
						 when  68  =>    DADOS_AUDIO <=  "0111110111000001";
						 when  69  =>    DADOS_AUDIO <=  "0111110100011001";
						 when  70  =>    DADOS_AUDIO <=  "0111110001011011";
						 when  71  =>    DADOS_AUDIO <=  "0111101110000111";
						 when  72  =>    DADOS_AUDIO <=  "0111101010011111";
						 when  73  =>    DADOS_AUDIO <=  "0111100110100001";
						 when  74  =>    DADOS_AUDIO <=  "0111100010001111";
						 when  75  =>    DADOS_AUDIO <=  "0111011101101000";
						 when  76  =>    DADOS_AUDIO <=  "0111011000101101";
						 when  77  =>    DADOS_AUDIO <=  "0111010011011101";
						 when  78  =>    DADOS_AUDIO <=  "0111001101111010";
						 when  79  =>    DADOS_AUDIO <=  "0111001000000010";
						 when  80  =>    DADOS_AUDIO <=  "0111000001111000";
						 when  81  =>    DADOS_AUDIO <=  "0110111011011001";
						 when  82  =>    DADOS_AUDIO <=  "0110110100101000";
						 when  83  =>    DADOS_AUDIO <=  "0110101101100101";
						 when  84  =>    DADOS_AUDIO <=  "0110100110001110";
						 when  85  =>    DADOS_AUDIO <=  "0110011110100110";
						 when  86  =>    DADOS_AUDIO <=  "0110010110101100";
						 when  87  =>    DADOS_AUDIO <=  "0110001110100001";
						 when  88  =>    DADOS_AUDIO <=  "0110000110000101";
						 when  89  =>    DADOS_AUDIO <=  "0101111101010111";
						 when  90  =>    DADOS_AUDIO <=  "0101110100011010";
						 when  91  =>    DADOS_AUDIO <=  "0101101011001101";
						 when  92  =>    DADOS_AUDIO <=  "0101100001110000";
						 when  93  =>    DADOS_AUDIO <=  "0101011000000100";
						 when  94  =>    DADOS_AUDIO <=  "0101001110001001";
						 when  95  =>    DADOS_AUDIO <=  "0101000100000000";
						 when  96  =>    DADOS_AUDIO <=  "0100111001101001";
						 when  97  =>    DADOS_AUDIO <=  "0100101111000101";
						 when  98  =>    DADOS_AUDIO <=  "0100100100010100";
						 when  99  =>    DADOS_AUDIO <=  "0100011001010110";
						 when  100  =>    DADOS_AUDIO <=  "0100001110001100";
						 when  101  =>    DADOS_AUDIO <=  "0100000010110111";
						 when  102  =>    DADOS_AUDIO <=  "0011110111010110";
						 when  103  =>    DADOS_AUDIO <=  "0011101011101011";
						 when  104  =>    DADOS_AUDIO <=  "0011011111110110";
						 when  105  =>    DADOS_AUDIO <=  "0011010011110111";
						 when  106  =>    DADOS_AUDIO <=  "0011000111101111";
						 when  107  =>    DADOS_AUDIO <=  "0010111011011111";
						 when  108  =>    DADOS_AUDIO <=  "0010101111000111";
						 when  109  =>    DADOS_AUDIO <=  "0010100010100111";
						 when  110  =>    DADOS_AUDIO <=  "0010010110000000";
						 when  111  =>    DADOS_AUDIO <=  "0010001001010011";
						 when  112  =>    DADOS_AUDIO <=  "0001111100100000";
						 when  113  =>    DADOS_AUDIO <=  "0001101111100111";
						 when  114  =>    DADOS_AUDIO <=  "0001100010101010";
						 when  115  =>    DADOS_AUDIO <=  "0001010101101001";
						 when  116  =>    DADOS_AUDIO <=  "0001001000100100";
						 when  117  =>    DADOS_AUDIO <=  "0000111011011100";
						 when  118  =>    DADOS_AUDIO <=  "0000101110010001";
						 when  119  =>    DADOS_AUDIO <=  "0000100001000100";
						 when  120  =>    DADOS_AUDIO <=  "0000010011110110";
						 when  121  =>    DADOS_AUDIO <=  "0000000110100111";
						 when  122  =>    DADOS_AUDIO <=  "1111111001011001";
						 when  123  =>    DADOS_AUDIO <=  "1111101100001010";
						 when  124  =>    DADOS_AUDIO <=  "1111011110111100";
						 when  125  =>    DADOS_AUDIO <=  "1111010001101111";
						 when  126  =>    DADOS_AUDIO <=  "1111000100100100";
						 when  127  =>    DADOS_AUDIO <=  "1110110111011100";
						 when  128  =>    DADOS_AUDIO <=  "1110101010010111";
						 when  129  =>    DADOS_AUDIO <=  "1110011101010110";
						 when  130  =>    DADOS_AUDIO <=  "1110010000011001";
						 when  131  =>    DADOS_AUDIO <=  "1110000011100000";
						 when  132  =>    DADOS_AUDIO <=  "1101110110101101";
						 when  133  =>    DADOS_AUDIO <=  "1101101010000000";
						 when  134  =>    DADOS_AUDIO <=  "1101011101011001";
						 when  135  =>    DADOS_AUDIO <=  "1101010000111001";
						 when  136  =>    DADOS_AUDIO <=  "1101000100100001";
						 when  137  =>    DADOS_AUDIO <=  "1100111000010001";
						 when  138  =>    DADOS_AUDIO <=  "1100101100001001";
						 when  139  =>    DADOS_AUDIO <=  "1100100000001010";
						 when  140  =>    DADOS_AUDIO <=  "1100010100010101";
						 when  141  =>    DADOS_AUDIO <=  "1100001000101010";
						 when  142  =>    DADOS_AUDIO <=  "1011111101001001";
						 when  143  =>    DADOS_AUDIO <=  "1011110001110100";
						 when  144  =>    DADOS_AUDIO <=  "1011100110101010";
						 when  145  =>    DADOS_AUDIO <=  "1011011011101100";
						 when  146  =>    DADOS_AUDIO <=  "1011010000111011";
						 when  147  =>    DADOS_AUDIO <=  "1011000110010111";
						 when  148  =>    DADOS_AUDIO <=  "1010111100000000";
						 when  149  =>    DADOS_AUDIO <=  "1010110001110111";
						 when  150  =>    DADOS_AUDIO <=  "1010100111111100";
						 when  151  =>    DADOS_AUDIO <=  "1010011110010000";
						 when  152  =>    DADOS_AUDIO <=  "1010010100110011";
						 when  153  =>    DADOS_AUDIO <=  "1010001011100110";
						 when  154  =>    DADOS_AUDIO <=  "1010000010101001";
						 when  155  =>    DADOS_AUDIO <=  "1001111001111011";
						 when  156  =>    DADOS_AUDIO <=  "1001110001011111";
						 when  157  =>    DADOS_AUDIO <=  "1001101001010100";
						 when  158  =>    DADOS_AUDIO <=  "1001100001011010";
						 when  159  =>    DADOS_AUDIO <=  "1001011001110010";
						 when  160  =>    DADOS_AUDIO <=  "1001010010011011";
						 when  161  =>    DADOS_AUDIO <=  "1001001011011000";
						 when  162  =>    DADOS_AUDIO <=  "1001000100100111";
						 when  163  =>    DADOS_AUDIO <=  "1000111110001000";
						 when  164  =>    DADOS_AUDIO <=  "1000110111111110";
						 when  165  =>    DADOS_AUDIO <=  "1000110010000110";
						 when  166  =>    DADOS_AUDIO <=  "1000101100100011";
						 when  167  =>    DADOS_AUDIO <=  "1000100111010011";
						 when  168  =>    DADOS_AUDIO <=  "1000100010011000";
						 when  169  =>    DADOS_AUDIO <=  "1000011101110001";
						 when  170  =>    DADOS_AUDIO <=  "1000011001011111";
						 when  171  =>    DADOS_AUDIO <=  "1000010101100001";
						 when  172  =>    DADOS_AUDIO <=  "1000010001111001";
						 when  173  =>    DADOS_AUDIO <=  "1000001110100101";
						 when  174  =>    DADOS_AUDIO <=  "1000001011100111";
						 when  175  =>    DADOS_AUDIO <=  "1000001000111111";
						 when  176  =>    DADOS_AUDIO <=  "1000000110101011";
						 when  177  =>    DADOS_AUDIO <=  "1000000100101110";
						 when  178  =>    DADOS_AUDIO <=  "1000000011000110";
						 when  179  =>    DADOS_AUDIO <=  "1000000001110100";
						 when  180  =>    DADOS_AUDIO <=  "1000000000111000";
						 when  181  =>    DADOS_AUDIO <=  "1000000000010010";
						 when  182  =>    DADOS_AUDIO <=  "1000000000000001";
						 when  183  =>    DADOS_AUDIO <=  "1000000000000111";
						 when  184  =>    DADOS_AUDIO <=  "1000000000100010";
						 when  185  =>    DADOS_AUDIO <=  "1000000001010011";
						 when  186  =>    DADOS_AUDIO <=  "1000000010011010";
						 when  187  =>    DADOS_AUDIO <=  "1000000011110111";
						 when  188  =>    DADOS_AUDIO <=  "1000000101101010";
						 when  189  =>    DADOS_AUDIO <=  "1000000111110010";
						 when  190  =>    DADOS_AUDIO <=  "1000001010010000";
						 when  191  =>    DADOS_AUDIO <=  "1000001101000100";
						 when  192  =>    DADOS_AUDIO <=  "1000010000001100";
						 when  193  =>    DADOS_AUDIO <=  "1000010011101010";
						 when  194  =>    DADOS_AUDIO <=  "1000010111011101";
						 when  195  =>    DADOS_AUDIO <=  "1000011011100101";
						 when  196  =>    DADOS_AUDIO <=  "1000100000000010";
						 when  197  =>    DADOS_AUDIO <=  "1000100100110011";
						 when  198  =>    DADOS_AUDIO <=  "1000101001111000";
						 when  199  =>    DADOS_AUDIO <=  "1000101111010010";
						 when  200  =>    DADOS_AUDIO <=  "1000110100111111";
						 when  201  =>    DADOS_AUDIO <=  "1000111011000001";
						 when  202  =>    DADOS_AUDIO <=  "1001000001010101";
						 when  203  =>    DADOS_AUDIO <=  "1001000111111101";
						 when  204  =>    DADOS_AUDIO <=  "1001001110110111";
						 when  205  =>    DADOS_AUDIO <=  "1001010110000100";
						 when  206  =>    DADOS_AUDIO <=  "1001011101100011";
						 when  207  =>    DADOS_AUDIO <=  "1001100101010101";
						 when  208  =>    DADOS_AUDIO <=  "1001101101010111";
						 when  209  =>    DADOS_AUDIO <=  "1001110101101011";
						 when  210  =>    DADOS_AUDIO <=  "1001111110010000";
						 when  211  =>    DADOS_AUDIO <=  "1010000111000101";
						 when  212  =>    DADOS_AUDIO <=  "1010010000001011";
						 when  213  =>    DADOS_AUDIO <=  "1010011001100000";
						 when  214  =>    DADOS_AUDIO <=  "1010100011000100";
						 when  215  =>    DADOS_AUDIO <=  "1010101100111000";
						 when  216  =>    DADOS_AUDIO <=  "1010110110111010";
						 when  217  =>    DADOS_AUDIO <=  "1011000001001010";
						 when  218  =>    DADOS_AUDIO <=  "1011001011100111";
						 when  219  =>    DADOS_AUDIO <=  "1011010110010010";
						 when  220  =>    DADOS_AUDIO <=  "1011100001001010";
						 when  221  =>    DADOS_AUDIO <=  "1011101100001110";
						 when  222  =>    DADOS_AUDIO <=  "1011110111011101";
						 when  223  =>    DADOS_AUDIO <=  "1100000010111000";
						 when  224  =>    DADOS_AUDIO <=  "1100001110011110";
						 when  225  =>    DADOS_AUDIO <=  "1100011010001110";
						 when  226  =>    DADOS_AUDIO <=  "1100100110001000";
						 when  227  =>    DADOS_AUDIO <=  "1100110010001100";
						 when  228  =>    DADOS_AUDIO <=  "1100111110011000";
						 when  229  =>    DADOS_AUDIO <=  "1101001010101100";
						 when  230  =>    DADOS_AUDIO <=  "1101010111001000";
						 when  231  =>    DADOS_AUDIO <=  "1101100011101100";
						 when  232  =>    DADOS_AUDIO <=  "1101110000010110";
						 when  233  =>    DADOS_AUDIO <=  "1101111101000110";
						 when  234  =>    DADOS_AUDIO <=  "1110001001111100";
						 when  235  =>    DADOS_AUDIO <=  "1110010110110111";
						 when  236  =>    DADOS_AUDIO <=  "1110100011110110";
						 when  237  =>    DADOS_AUDIO <=  "1110110000111001";
						 when  238  =>    DADOS_AUDIO <=  "1110111110000000";
						 when  239  =>    DADOS_AUDIO <=  "1111001011001001";
						 when  240  =>    DADOS_AUDIO <=  "1111011000010101";
						 when  241  =>    DADOS_AUDIO <=  "1111100101100011";
						 when  242  =>    DADOS_AUDIO <=  "1111110010110001";
						 when  243  =>    DADOS_AUDIO <=  "0000000000000000";
						 when others =>	DADOS_AUDIO <=  "0000000000000000";
					end case;
				when 9 =>
					n_pontos <= 231;
					reset <= '0';
					case aux_dados is
					    when  0  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  1  =>    DADOS_AUDIO <=  "0000001101111111";
						 when  2  =>    DADOS_AUDIO <=  "0000011011111101";
						 when  3  =>    DADOS_AUDIO <=  "0000101001111010";
						 when  4  =>    DADOS_AUDIO <=  "0000110111110101";
						 when  5  =>    DADOS_AUDIO <=  "0001000101101101";
						 when  6  =>    DADOS_AUDIO <=  "0001010011100010";
						 when  7  =>    DADOS_AUDIO <=  "0001100001010100";
						 when  8  =>    DADOS_AUDIO <=  "0001101111000000";
						 when  9  =>    DADOS_AUDIO <=  "0001111100100111";
						 when  10  =>    DADOS_AUDIO <=  "0010001010001000";
						 when  11  =>    DADOS_AUDIO <=  "0010010111100011";
						 when  12  =>    DADOS_AUDIO <=  "0010100100110110";
						 when  13  =>    DADOS_AUDIO <=  "0010110010000010";
						 when  14  =>    DADOS_AUDIO <=  "0010111111000100";
						 when  15  =>    DADOS_AUDIO <=  "0011001011111110";
						 when  16  =>    DADOS_AUDIO <=  "0011011000101110";
						 when  17  =>    DADOS_AUDIO <=  "0011100101010100";
						 when  18  =>    DADOS_AUDIO <=  "0011110001101111";
						 when  19  =>    DADOS_AUDIO <=  "0011111101111110";
						 when  20  =>    DADOS_AUDIO <=  "0100001010000001";
						 when  21  =>    DADOS_AUDIO <=  "0100010101111000";
						 when  22  =>    DADOS_AUDIO <=  "0100100001100001";
						 when  23  =>    DADOS_AUDIO <=  "0100101100111100";
						 when  24  =>    DADOS_AUDIO <=  "0100111000001001";
						 when  25  =>    DADOS_AUDIO <=  "0101000011000111";
						 when  26  =>    DADOS_AUDIO <=  "0101001101110110";
						 when  27  =>    DADOS_AUDIO <=  "0101011000010100";
						 when  28  =>    DADOS_AUDIO <=  "0101100010100010";
						 when  29  =>    DADOS_AUDIO <=  "0101101100100000";
						 when  30  =>    DADOS_AUDIO <=  "0101110110001100";
						 when  31  =>    DADOS_AUDIO <=  "0101111111100110";
						 when  32  =>    DADOS_AUDIO <=  "0110001000101101";
						 when  33  =>    DADOS_AUDIO <=  "0110010001100010";
						 when  34  =>    DADOS_AUDIO <=  "0110011010000100";
						 when  35  =>    DADOS_AUDIO <=  "0110100010010010";
						 when  36  =>    DADOS_AUDIO <=  "0110101010001100";
						 when  37  =>    DADOS_AUDIO <=  "0110110001110010";
						 when  38  =>    DADOS_AUDIO <=  "0110111001000011";
						 when  39  =>    DADOS_AUDIO <=  "0110111111111111";
						 when  40  =>    DADOS_AUDIO <=  "0111000110100110";
						 when  41  =>    DADOS_AUDIO <=  "0111001100110111";
						 when  42  =>    DADOS_AUDIO <=  "0111010010110010";
						 when  43  =>    DADOS_AUDIO <=  "0111011000010110";
						 when  44  =>    DADOS_AUDIO <=  "0111011101100100";
						 when  45  =>    DADOS_AUDIO <=  "0111100010011100";
						 when  46  =>    DADOS_AUDIO <=  "0111100110111100";
						 when  47  =>    DADOS_AUDIO <=  "0111101011000101";
						 when  48  =>    DADOS_AUDIO <=  "0111101110110110";
						 when  49  =>    DADOS_AUDIO <=  "0111110010010000";
						 when  50  =>    DADOS_AUDIO <=  "0111110101010010";
						 when  51  =>    DADOS_AUDIO <=  "0111110111111100";
						 when  52  =>    DADOS_AUDIO <=  "0111111010001110";
						 when  53  =>    DADOS_AUDIO <=  "0111111100001000";
						 when  54  =>    DADOS_AUDIO <=  "0111111101101010";
						 when  55  =>    DADOS_AUDIO <=  "0111111110110011";
						 when  56  =>    DADOS_AUDIO <=  "0111111111100100";
						 when  57  =>    DADOS_AUDIO <=  "0111111111111100";
						 when  58  =>    DADOS_AUDIO <=  "0111111111111100";
						 when  59  =>    DADOS_AUDIO <=  "0111111111100100";
						 when  60  =>    DADOS_AUDIO <=  "0111111110110011";
						 when  61  =>    DADOS_AUDIO <=  "0111111101101010";
						 when  62  =>    DADOS_AUDIO <=  "0111111100001000";
						 when  63  =>    DADOS_AUDIO <=  "0111111010001110";
						 when  64  =>    DADOS_AUDIO <=  "0111110111111100";
						 when  65  =>    DADOS_AUDIO <=  "0111110101010010";
						 when  66  =>    DADOS_AUDIO <=  "0111110010010000";
						 when  67  =>    DADOS_AUDIO <=  "0111101110110110";
						 when  68  =>    DADOS_AUDIO <=  "0111101011000101";
						 when  69  =>    DADOS_AUDIO <=  "0111100110111100";
						 when  70  =>    DADOS_AUDIO <=  "0111100010011100";
						 when  71  =>    DADOS_AUDIO <=  "0111011101100100";
						 when  72  =>    DADOS_AUDIO <=  "0111011000010110";
						 when  73  =>    DADOS_AUDIO <=  "0111010010110010";
						 when  74  =>    DADOS_AUDIO <=  "0111001100110111";
						 when  75  =>    DADOS_AUDIO <=  "0111000110100110";
						 when  76  =>    DADOS_AUDIO <=  "0110111111111111";
						 when  77  =>    DADOS_AUDIO <=  "0110111001000011";
						 when  78  =>    DADOS_AUDIO <=  "0110110001110010";
						 when  79  =>    DADOS_AUDIO <=  "0110101010001100";
						 when  80  =>    DADOS_AUDIO <=  "0110100010010010";
						 when  81  =>    DADOS_AUDIO <=  "0110011010000100";
						 when  82  =>    DADOS_AUDIO <=  "0110010001100010";
						 when  83  =>    DADOS_AUDIO <=  "0110001000101101";
						 when  84  =>    DADOS_AUDIO <=  "0101111111100110";
						 when  85  =>    DADOS_AUDIO <=  "0101110110001100";
						 when  86  =>    DADOS_AUDIO <=  "0101101100100000";
						 when  87  =>    DADOS_AUDIO <=  "0101100010100010";
						 when  88  =>    DADOS_AUDIO <=  "0101011000010100";
						 when  89  =>    DADOS_AUDIO <=  "0101001101110110";
						 when  90  =>    DADOS_AUDIO <=  "0101000011000111";
						 when  91  =>    DADOS_AUDIO <=  "0100111000001001";
						 when  92  =>    DADOS_AUDIO <=  "0100101100111100";
						 when  93  =>    DADOS_AUDIO <=  "0100100001100001";
						 when  94  =>    DADOS_AUDIO <=  "0100010101111000";
						 when  95  =>    DADOS_AUDIO <=  "0100001010000001";
						 when  96  =>    DADOS_AUDIO <=  "0011111101111110";
						 when  97  =>    DADOS_AUDIO <=  "0011110001101111";
						 when  98  =>    DADOS_AUDIO <=  "0011100101010100";
						 when  99  =>    DADOS_AUDIO <=  "0011011000101110";
						 when  100  =>    DADOS_AUDIO <=  "0011001011111110";
						 when  101  =>    DADOS_AUDIO <=  "0010111111000100";
						 when  102  =>    DADOS_AUDIO <=  "0010110010000010";
						 when  103  =>    DADOS_AUDIO <=  "0010100100110110";
						 when  104  =>    DADOS_AUDIO <=  "0010010111100011";
						 when  105  =>    DADOS_AUDIO <=  "0010001010001000";
						 when  106  =>    DADOS_AUDIO <=  "0001111100100111";
						 when  107  =>    DADOS_AUDIO <=  "0001101111000000";
						 when  108  =>    DADOS_AUDIO <=  "0001100001010100";
						 when  109  =>    DADOS_AUDIO <=  "0001010011100010";
						 when  110  =>    DADOS_AUDIO <=  "0001000101101101";
						 when  111  =>    DADOS_AUDIO <=  "0000110111110101";
						 when  112  =>    DADOS_AUDIO <=  "0000101001111010";
						 when  113  =>    DADOS_AUDIO <=  "0000011011111101";
						 when  114  =>    DADOS_AUDIO <=  "0000001101111111";
						 when  115  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  116  =>    DADOS_AUDIO <=  "1111110010000001";
						 when  117  =>    DADOS_AUDIO <=  "1111100100000011";
						 when  118  =>    DADOS_AUDIO <=  "1111010110000110";
						 when  119  =>    DADOS_AUDIO <=  "1111001000001011";
						 when  120  =>    DADOS_AUDIO <=  "1110111010010011";
						 when  121  =>    DADOS_AUDIO <=  "1110101100011110";
						 when  122  =>    DADOS_AUDIO <=  "1110011110101100";
						 when  123  =>    DADOS_AUDIO <=  "1110010001000000";
						 when  124  =>    DADOS_AUDIO <=  "1110000011011001";
						 when  125  =>    DADOS_AUDIO <=  "1101110101111000";
						 when  126  =>    DADOS_AUDIO <=  "1101101000011101";
						 when  127  =>    DADOS_AUDIO <=  "1101011011001010";
						 when  128  =>    DADOS_AUDIO <=  "1101001101111110";
						 when  129  =>    DADOS_AUDIO <=  "1101000000111100";
						 when  130  =>    DADOS_AUDIO <=  "1100110100000010";
						 when  131  =>    DADOS_AUDIO <=  "1100100111010010";
						 when  132  =>    DADOS_AUDIO <=  "1100011010101100";
						 when  133  =>    DADOS_AUDIO <=  "1100001110010001";
						 when  134  =>    DADOS_AUDIO <=  "1100000010000010";
						 when  135  =>    DADOS_AUDIO <=  "1011110101111111";
						 when  136  =>    DADOS_AUDIO <=  "1011101010001000";
						 when  137  =>    DADOS_AUDIO <=  "1011011110011111";
						 when  138  =>    DADOS_AUDIO <=  "1011010011000100";
						 when  139  =>    DADOS_AUDIO <=  "1011000111110111";
						 when  140  =>    DADOS_AUDIO <=  "1010111100111001";
						 when  141  =>    DADOS_AUDIO <=  "1010110010001010";
						 when  142  =>    DADOS_AUDIO <=  "1010100111101100";
						 when  143  =>    DADOS_AUDIO <=  "1010011101011110";
						 when  144  =>    DADOS_AUDIO <=  "1010010011100000";
						 when  145  =>    DADOS_AUDIO <=  "1010001001110100";
						 when  146  =>    DADOS_AUDIO <=  "1010000000011010";
						 when  147  =>    DADOS_AUDIO <=  "1001110111010011";
						 when  148  =>    DADOS_AUDIO <=  "1001101110011110";
						 when  149  =>    DADOS_AUDIO <=  "1001100101111100";
						 when  150  =>    DADOS_AUDIO <=  "1001011101101110";
						 when  151  =>    DADOS_AUDIO <=  "1001010101110100";
						 when  152  =>    DADOS_AUDIO <=  "1001001110001110";
						 when  153  =>    DADOS_AUDIO <=  "1001000110111101";
						 when  154  =>    DADOS_AUDIO <=  "1001000000000001";
						 when  155  =>    DADOS_AUDIO <=  "1000111001011010";
						 when  156  =>    DADOS_AUDIO <=  "1000110011001001";
						 when  157  =>    DADOS_AUDIO <=  "1000101101001110";
						 when  158  =>    DADOS_AUDIO <=  "1000100111101010";
						 when  159  =>    DADOS_AUDIO <=  "1000100010011100";
						 when  160  =>    DADOS_AUDIO <=  "1000011101100100";
						 when  161  =>    DADOS_AUDIO <=  "1000011001000100";
						 when  162  =>    DADOS_AUDIO <=  "1000010100111011";
						 when  163  =>    DADOS_AUDIO <=  "1000010001001010";
						 when  164  =>    DADOS_AUDIO <=  "1000001101110000";
						 when  165  =>    DADOS_AUDIO <=  "1000001010101110";
						 when  166  =>    DADOS_AUDIO <=  "1000001000000100";
						 when  167  =>    DADOS_AUDIO <=  "1000000101110010";
						 when  168  =>    DADOS_AUDIO <=  "1000000011111000";
						 when  169  =>    DADOS_AUDIO <=  "1000000010010110";
						 when  170  =>    DADOS_AUDIO <=  "1000000001001101";
						 when  171  =>    DADOS_AUDIO <=  "1000000000011100";
						 when  172  =>    DADOS_AUDIO <=  "1000000000000100";
						 when  173  =>    DADOS_AUDIO <=  "1000000000000100";
						 when  174  =>    DADOS_AUDIO <=  "1000000000011100";
						 when  175  =>    DADOS_AUDIO <=  "1000000001001101";
						 when  176  =>    DADOS_AUDIO <=  "1000000010010110";
						 when  177  =>    DADOS_AUDIO <=  "1000000011111000";
						 when  178  =>    DADOS_AUDIO <=  "1000000101110010";
						 when  179  =>    DADOS_AUDIO <=  "1000001000000100";
						 when  180  =>    DADOS_AUDIO <=  "1000001010101110";
						 when  181  =>    DADOS_AUDIO <=  "1000001101110000";
						 when  182  =>    DADOS_AUDIO <=  "1000010001001010";
						 when  183  =>    DADOS_AUDIO <=  "1000010100111011";
						 when  184  =>    DADOS_AUDIO <=  "1000011001000100";
						 when  185  =>    DADOS_AUDIO <=  "1000011101100100";
						 when  186  =>    DADOS_AUDIO <=  "1000100010011100";
						 when  187  =>    DADOS_AUDIO <=  "1000100111101010";
						 when  188  =>    DADOS_AUDIO <=  "1000101101001110";
						 when  189  =>    DADOS_AUDIO <=  "1000110011001001";
						 when  190  =>    DADOS_AUDIO <=  "1000111001011010";
						 when  191  =>    DADOS_AUDIO <=  "1001000000000001";
						 when  192  =>    DADOS_AUDIO <=  "1001000110111101";
						 when  193  =>    DADOS_AUDIO <=  "1001001110001110";
						 when  194  =>    DADOS_AUDIO <=  "1001010101110100";
						 when  195  =>    DADOS_AUDIO <=  "1001011101101110";
						 when  196  =>    DADOS_AUDIO <=  "1001100101111100";
						 when  197  =>    DADOS_AUDIO <=  "1001101110011110";
						 when  198  =>    DADOS_AUDIO <=  "1001110111010011";
						 when  199  =>    DADOS_AUDIO <=  "1010000000011010";
						 when  200  =>    DADOS_AUDIO <=  "1010001001110100";
						 when  201  =>    DADOS_AUDIO <=  "1010010011100000";
						 when  202  =>    DADOS_AUDIO <=  "1010011101011110";
						 when  203  =>    DADOS_AUDIO <=  "1010100111101100";
						 when  204  =>    DADOS_AUDIO <=  "1010110010001010";
						 when  205  =>    DADOS_AUDIO <=  "1010111100111001";
						 when  206  =>    DADOS_AUDIO <=  "1011000111110111";
						 when  207  =>    DADOS_AUDIO <=  "1011010011000100";
						 when  208  =>    DADOS_AUDIO <=  "1011011110011111";
						 when  209  =>    DADOS_AUDIO <=  "1011101010001000";
						 when  210  =>    DADOS_AUDIO <=  "1011110101111111";
						 when  211  =>    DADOS_AUDIO <=  "1100000010000010";
						 when  212  =>    DADOS_AUDIO <=  "1100001110010001";
						 when  213  =>    DADOS_AUDIO <=  "1100011010101100";
						 when  214  =>    DADOS_AUDIO <=  "1100100111010010";
						 when  215  =>    DADOS_AUDIO <=  "1100110100000010";
						 when  216  =>    DADOS_AUDIO <=  "1101000000111100";
						 when  217  =>    DADOS_AUDIO <=  "1101001101111110";
						 when  218  =>    DADOS_AUDIO <=  "1101011011001010";
						 when  219  =>    DADOS_AUDIO <=  "1101101000011101";
						 when  220  =>    DADOS_AUDIO <=  "1101110101111000";
						 when  221  =>    DADOS_AUDIO <=  "1110000011011001";
						 when  222  =>    DADOS_AUDIO <=  "1110010001000000";
						 when  223  =>    DADOS_AUDIO <=  "1110011110101100";
						 when  224  =>    DADOS_AUDIO <=  "1110101100011110";
						 when  225  =>    DADOS_AUDIO <=  "1110111010010011";
						 when  226  =>    DADOS_AUDIO <=  "1111001000001011";
						 when  227  =>    DADOS_AUDIO <=  "1111010110000110";
						 when  228  =>    DADOS_AUDIO <=  "1111100100000011";
						 when  229  =>    DADOS_AUDIO <=  "1111110010000001";
						 when  230  =>    DADOS_AUDIO <=  "0000000000000000";
						 when others =>	DADOS_AUDIO <=  "0000000000000000";
					end case;
				when 10 =>
					n_pontos <= 218;
					reset <= '0';
					case aux_dados is
					    when  0  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  1  =>    DADOS_AUDIO <=  "0000001110110100";
						 when  2  =>    DADOS_AUDIO <=  "0000011101101000";
						 when  3  =>    DADOS_AUDIO <=  "0000101100011010";
						 when  4  =>    DADOS_AUDIO <=  "0000111011001010";
						 when  5  =>    DADOS_AUDIO <=  "0001001001110111";
						 when  6  =>    DADOS_AUDIO <=  "0001011000100000";
						 when  7  =>    DADOS_AUDIO <=  "0001100111000100";
						 when  8  =>    DADOS_AUDIO <=  "0001110101100010";
						 when  9  =>    DADOS_AUDIO <=  "0010000011111010";
						 when  10  =>    DADOS_AUDIO <=  "0010010010001011";
						 when  11  =>    DADOS_AUDIO <=  "0010100000010101";
						 when  12  =>    DADOS_AUDIO <=  "0010101110010101";
						 when  13  =>    DADOS_AUDIO <=  "0010111100001101";
						 when  14  =>    DADOS_AUDIO <=  "0011001001111010";
						 when  15  =>    DADOS_AUDIO <=  "0011010111011100";
						 when  16  =>    DADOS_AUDIO <=  "0011100100110011";
						 when  17  =>    DADOS_AUDIO <=  "0011110001111101";
						 when  18  =>    DADOS_AUDIO <=  "0011111110111011";
						 when  19  =>    DADOS_AUDIO <=  "0100001011101011";
						 when  20  =>    DADOS_AUDIO <=  "0100011000001100";
						 when  21  =>    DADOS_AUDIO <=  "0100100100011111";
						 when  22  =>    DADOS_AUDIO <=  "0100110000100010";
						 when  23  =>    DADOS_AUDIO <=  "0100111100010100";
						 when  24  =>    DADOS_AUDIO <=  "0101000111110101";
						 when  25  =>    DADOS_AUDIO <=  "0101010011000101";
						 when  26  =>    DADOS_AUDIO <=  "0101011110000011";
						 when  27  =>    DADOS_AUDIO <=  "0101101000101110";
						 when  28  =>    DADOS_AUDIO <=  "0101110011000110";
						 when  29  =>    DADOS_AUDIO <=  "0101111101001001";
						 when  30  =>    DADOS_AUDIO <=  "0110000110111000";
						 when  31  =>    DADOS_AUDIO <=  "0110010000010011";
						 when  32  =>    DADOS_AUDIO <=  "0110011001010111";
						 when  33  =>    DADOS_AUDIO <=  "0110100010000110";
						 when  34  =>    DADOS_AUDIO <=  "0110101010011110";
						 when  35  =>    DADOS_AUDIO <=  "0110110010100000";
						 when  36  =>    DADOS_AUDIO <=  "0110111010001010";
						 when  37  =>    DADOS_AUDIO <=  "0111000001011100";
						 when  38  =>    DADOS_AUDIO <=  "0111001000010111";
						 when  39  =>    DADOS_AUDIO <=  "0111001110111001";
						 when  40  =>    DADOS_AUDIO <=  "0111010101000010";
						 when  41  =>    DADOS_AUDIO <=  "0111011010110001";
						 when  42  =>    DADOS_AUDIO <=  "0111100000001000";
						 when  43  =>    DADOS_AUDIO <=  "0111100101000100";
						 when  44  =>    DADOS_AUDIO <=  "0111101001100111";
						 when  45  =>    DADOS_AUDIO <=  "0111101101101111";
						 when  46  =>    DADOS_AUDIO <=  "0111110001011101";
						 when  47  =>    DADOS_AUDIO <=  "0111110100110000";
						 when  48  =>    DADOS_AUDIO <=  "0111110111101000";
						 when  49  =>    DADOS_AUDIO <=  "0111111010000110";
						 when  50  =>    DADOS_AUDIO <=  "0111111100001000";
						 when  51  =>    DADOS_AUDIO <=  "0111111101101111";
						 when  52  =>    DADOS_AUDIO <=  "0111111110111010";
						 when  53  =>    DADOS_AUDIO <=  "0111111111101010";
						 when  54  =>    DADOS_AUDIO <=  "0111111111111111";
						 when  55  =>    DADOS_AUDIO <=  "0111111111111000";
						 when  56  =>    DADOS_AUDIO <=  "0111111111010101";
						 when  57  =>    DADOS_AUDIO <=  "0111111110011000";
						 when  58  =>    DADOS_AUDIO <=  "0111111100111111";
						 when  59  =>    DADOS_AUDIO <=  "0111111011001010";
						 when  60  =>    DADOS_AUDIO <=  "0111111000111010";
						 when  61  =>    DADOS_AUDIO <=  "0111110110010000";
						 when  62  =>    DADOS_AUDIO <=  "0111110011001010";
						 when  63  =>    DADOS_AUDIO <=  "0111101111101001";
						 when  64  =>    DADOS_AUDIO <=  "0111101011101110";
						 when  65  =>    DADOS_AUDIO <=  "0111100111011001";
						 when  66  =>    DADOS_AUDIO <=  "0111100010101001";
						 when  67  =>    DADOS_AUDIO <=  "0111011101100000";
						 when  68  =>    DADOS_AUDIO <=  "0111010111111101";
						 when  69  =>    DADOS_AUDIO <=  "0111010010000000";
						 when  70  =>    DADOS_AUDIO <=  "0111001011101011";
						 when  71  =>    DADOS_AUDIO <=  "0111000100111101";
						 when  72  =>    DADOS_AUDIO <=  "0110111101110110";
						 when  73  =>    DADOS_AUDIO <=  "0110110110011000";
						 when  74  =>    DADOS_AUDIO <=  "0110101110100010";
						 when  75  =>    DADOS_AUDIO <=  "0110100110010101";
						 when  76  =>    DADOS_AUDIO <=  "0110011101110001";
						 when  77  =>    DADOS_AUDIO <=  "0110010100111000";
						 when  78  =>    DADOS_AUDIO <=  "0110001011101000";
						 when  79  =>    DADOS_AUDIO <=  "0110000010000011";
						 when  80  =>    DADOS_AUDIO <=  "0101111000001010";
						 when  81  =>    DADOS_AUDIO <=  "0101101101111100";
						 when  82  =>    DADOS_AUDIO <=  "0101100011011011";
						 when  83  =>    DADOS_AUDIO <=  "0101011000100111";
						 when  84  =>    DADOS_AUDIO <=  "0101001101100000";
						 when  85  =>    DADOS_AUDIO <=  "0101000010000111";
						 when  86  =>    DADOS_AUDIO <=  "0100110110011101";
						 when  87  =>    DADOS_AUDIO <=  "0100101010100010";
						 when  88  =>    DADOS_AUDIO <=  "0100011110011000";
						 when  89  =>    DADOS_AUDIO <=  "0100010001111101";
						 when  90  =>    DADOS_AUDIO <=  "0100000101010101";
						 when  91  =>    DADOS_AUDIO <=  "0011111000011110";
						 when  92  =>    DADOS_AUDIO <=  "0011101011011010";
						 when  93  =>    DADOS_AUDIO <=  "0011011110001001";
						 when  94  =>    DADOS_AUDIO <=  "0011010000101100";
						 when  95  =>    DADOS_AUDIO <=  "0011000011000100";
						 when  96  =>    DADOS_AUDIO <=  "0010110101010010";
						 when  97  =>    DADOS_AUDIO <=  "0010100111010110";
						 when  98  =>    DADOS_AUDIO <=  "0010011001010001";
						 when  99  =>    DADOS_AUDIO <=  "0010001011000100";
						 when  100  =>    DADOS_AUDIO <=  "0001111100101111";
						 when  101  =>    DADOS_AUDIO <=  "0001101110010100";
						 when  102  =>    DADOS_AUDIO <=  "0001011111110010";
						 when  103  =>    DADOS_AUDIO <=  "0001010001001100";
						 when  104  =>    DADOS_AUDIO <=  "0001000010100001";
						 when  105  =>    DADOS_AUDIO <=  "0000110011110011";
						 when  106  =>    DADOS_AUDIO <=  "0000100101000001";
						 when  107  =>    DADOS_AUDIO <=  "0000010110001110";
						 when  108  =>    DADOS_AUDIO <=  "0000000111011010";
						 when  109  =>    DADOS_AUDIO <=  "1111111000100110";
						 when  110  =>    DADOS_AUDIO <=  "1111101001110010";
						 when  111  =>    DADOS_AUDIO <=  "1111011010111111";
						 when  112  =>    DADOS_AUDIO <=  "1111001100001101";
						 when  113  =>    DADOS_AUDIO <=  "1110111101011111";
						 when  114  =>    DADOS_AUDIO <=  "1110101110110100";
						 when  115  =>    DADOS_AUDIO <=  "1110100000001110";
						 when  116  =>    DADOS_AUDIO <=  "1110010001101100";
						 when  117  =>    DADOS_AUDIO <=  "1110000011010001";
						 when  118  =>    DADOS_AUDIO <=  "1101110100111100";
						 when  119  =>    DADOS_AUDIO <=  "1101100110101111";
						 when  120  =>    DADOS_AUDIO <=  "1101011000101010";
						 when  121  =>    DADOS_AUDIO <=  "1101001010101110";
						 when  122  =>    DADOS_AUDIO <=  "1100111100111100";
						 when  123  =>    DADOS_AUDIO <=  "1100101111010100";
						 when  124  =>    DADOS_AUDIO <=  "1100100001110111";
						 when  125  =>    DADOS_AUDIO <=  "1100010100100110";
						 when  126  =>    DADOS_AUDIO <=  "1100000111100010";
						 when  127  =>    DADOS_AUDIO <=  "1011111010101011";
						 when  128  =>    DADOS_AUDIO <=  "1011101110000011";
						 when  129  =>    DADOS_AUDIO <=  "1011100001101000";
						 when  130  =>    DADOS_AUDIO <=  "1011010101011110";
						 when  131  =>    DADOS_AUDIO <=  "1011001001100011";
						 when  132  =>    DADOS_AUDIO <=  "1010111101111001";
						 when  133  =>    DADOS_AUDIO <=  "1010110010100000";
						 when  134  =>    DADOS_AUDIO <=  "1010100111011001";
						 when  135  =>    DADOS_AUDIO <=  "1010011100100101";
						 when  136  =>    DADOS_AUDIO <=  "1010010010000100";
						 when  137  =>    DADOS_AUDIO <=  "1010000111110110";
						 when  138  =>    DADOS_AUDIO <=  "1001111101111101";
						 when  139  =>    DADOS_AUDIO <=  "1001110100011000";
						 when  140  =>    DADOS_AUDIO <=  "1001101011001000";
						 when  141  =>    DADOS_AUDIO <=  "1001100010001111";
						 when  142  =>    DADOS_AUDIO <=  "1001011001101011";
						 when  143  =>    DADOS_AUDIO <=  "1001010001011110";
						 when  144  =>    DADOS_AUDIO <=  "1001001001101000";
						 when  145  =>    DADOS_AUDIO <=  "1001000010001010";
						 when  146  =>    DADOS_AUDIO <=  "1000111011000011";
						 when  147  =>    DADOS_AUDIO <=  "1000110100010101";
						 when  148  =>    DADOS_AUDIO <=  "1000101110000000";
						 when  149  =>    DADOS_AUDIO <=  "1000101000000011";
						 when  150  =>    DADOS_AUDIO <=  "1000100010100000";
						 when  151  =>    DADOS_AUDIO <=  "1000011101010111";
						 when  152  =>    DADOS_AUDIO <=  "1000011000100111";
						 when  153  =>    DADOS_AUDIO <=  "1000010100010010";
						 when  154  =>    DADOS_AUDIO <=  "1000010000010111";
						 when  155  =>    DADOS_AUDIO <=  "1000001100110110";
						 when  156  =>    DADOS_AUDIO <=  "1000001001110000";
						 when  157  =>    DADOS_AUDIO <=  "1000000111000110";
						 when  158  =>    DADOS_AUDIO <=  "1000000100110110";
						 when  159  =>    DADOS_AUDIO <=  "1000000011000001";
						 when  160  =>    DADOS_AUDIO <=  "1000000001101000";
						 when  161  =>    DADOS_AUDIO <=  "1000000000101011";
						 when  162  =>    DADOS_AUDIO <=  "1000000000001000";
						 when  163  =>    DADOS_AUDIO <=  "1000000000000001";
						 when  164  =>    DADOS_AUDIO <=  "1000000000010110";
						 when  165  =>    DADOS_AUDIO <=  "1000000001000110";
						 when  166  =>    DADOS_AUDIO <=  "1000000010010001";
						 when  167  =>    DADOS_AUDIO <=  "1000000011111000";
						 when  168  =>    DADOS_AUDIO <=  "1000000101111010";
						 when  169  =>    DADOS_AUDIO <=  "1000001000011000";
						 when  170  =>    DADOS_AUDIO <=  "1000001011010000";
						 when  171  =>    DADOS_AUDIO <=  "1000001110100011";
						 when  172  =>    DADOS_AUDIO <=  "1000010010010001";
						 when  173  =>    DADOS_AUDIO <=  "1000010110011001";
						 when  174  =>    DADOS_AUDIO <=  "1000011010111100";
						 when  175  =>    DADOS_AUDIO <=  "1000011111111000";
						 when  176  =>    DADOS_AUDIO <=  "1000100101001111";
						 when  177  =>    DADOS_AUDIO <=  "1000101010111110";
						 when  178  =>    DADOS_AUDIO <=  "1000110001000111";
						 when  179  =>    DADOS_AUDIO <=  "1000110111101001";
						 when  180  =>    DADOS_AUDIO <=  "1000111110100100";
						 when  181  =>    DADOS_AUDIO <=  "1001000101110110";
						 when  182  =>    DADOS_AUDIO <=  "1001001101100000";
						 when  183  =>    DADOS_AUDIO <=  "1001010101100010";
						 when  184  =>    DADOS_AUDIO <=  "1001011101111010";
						 when  185  =>    DADOS_AUDIO <=  "1001100110101001";
						 when  186  =>    DADOS_AUDIO <=  "1001101111101101";
						 when  187  =>    DADOS_AUDIO <=  "1001111001001000";
						 when  188  =>    DADOS_AUDIO <=  "1010000010110111";
						 when  189  =>    DADOS_AUDIO <=  "1010001100111010";
						 when  190  =>    DADOS_AUDIO <=  "1010010111010010";
						 when  191  =>    DADOS_AUDIO <=  "1010100001111101";
						 when  192  =>    DADOS_AUDIO <=  "1010101100111011";
						 when  193  =>    DADOS_AUDIO <=  "1010111000001011";
						 when  194  =>    DADOS_AUDIO <=  "1011000011101100";
						 when  195  =>    DADOS_AUDIO <=  "1011001111011110";
						 when  196  =>    DADOS_AUDIO <=  "1011011011100001";
						 when  197  =>    DADOS_AUDIO <=  "1011100111110100";
						 when  198  =>    DADOS_AUDIO <=  "1011110100010101";
						 when  199  =>    DADOS_AUDIO <=  "1100000001000101";
						 when  200  =>    DADOS_AUDIO <=  "1100001110000011";
						 when  201  =>    DADOS_AUDIO <=  "1100011011001101";
						 when  202  =>    DADOS_AUDIO <=  "1100101000100100";
						 when  203  =>    DADOS_AUDIO <=  "1100110110000110";
						 when  204  =>    DADOS_AUDIO <=  "1101000011110011";
						 when  205  =>    DADOS_AUDIO <=  "1101010001101011";
						 when  206  =>    DADOS_AUDIO <=  "1101011111101011";
						 when  207  =>    DADOS_AUDIO <=  "1101101101110101";
						 when  208  =>    DADOS_AUDIO <=  "1101111100000110";
						 when  209  =>    DADOS_AUDIO <=  "1110001010011110";
						 when  210  =>    DADOS_AUDIO <=  "1110011000111100";
						 when  211  =>    DADOS_AUDIO <=  "1110100111100000";
						 when  212  =>    DADOS_AUDIO <=  "1110110110001001";
						 when  213  =>    DADOS_AUDIO <=  "1111000100110110";
						 when  214  =>    DADOS_AUDIO <=  "1111010011100110";
						 when  215  =>    DADOS_AUDIO <=  "1111100010011000";
						 when  216  =>    DADOS_AUDIO <=  "1111110001001100";
						 when  217  =>    DADOS_AUDIO <=  "0000000000000000";
						 when others =>	DADOS_AUDIO <=  "0000000000000000";
					end case;
				when 11 =>
					n_pontos <= 206;
					reset <= '0';
					case aux_dados is
					    when  0  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  1  =>    DADOS_AUDIO <=  "0000001111101100";
						 when  2  =>    DADOS_AUDIO <=  "0000011111010111";
						 when  3  =>    DADOS_AUDIO <=  "0000101111000000";
						 when  4  =>    DADOS_AUDIO <=  "0000111110100111";
						 when  5  =>    DADOS_AUDIO <=  "0001001110001010";
						 when  6  =>    DADOS_AUDIO <=  "0001011101101000";
						 when  7  =>    DADOS_AUDIO <=  "0001101101000000";
						 when  8  =>    DADOS_AUDIO <=  "0001111100010010";
						 when  9  =>    DADOS_AUDIO <=  "0010001011011100";
						 when  10  =>    DADOS_AUDIO <=  "0010011010011110";
						 when  11  =>    DADOS_AUDIO <=  "0010101001010111";
						 when  12  =>    DADOS_AUDIO <=  "0010111000000110";
						 when  13  =>    DADOS_AUDIO <=  "0011000110101001";
						 when  14  =>    DADOS_AUDIO <=  "0011010101000001";
						 when  15  =>    DADOS_AUDIO <=  "0011100011001011";
						 when  16  =>    DADOS_AUDIO <=  "0011110001001000";
						 when  17  =>    DADOS_AUDIO <=  "0011111110110111";
						 when  18  =>    DADOS_AUDIO <=  "0100001100010110";
						 when  19  =>    DADOS_AUDIO <=  "0100011001100101";
						 when  20  =>    DADOS_AUDIO <=  "0100100110100100";
						 when  21  =>    DADOS_AUDIO <=  "0100110011010000";
						 when  22  =>    DADOS_AUDIO <=  "0100111111101010";
						 when  23  =>    DADOS_AUDIO <=  "0101001011110001";
						 when  24  =>    DADOS_AUDIO <=  "0101010111100100";
						 when  25  =>    DADOS_AUDIO <=  "0101100011000010";
						 when  26  =>    DADOS_AUDIO <=  "0101101110001011";
						 when  27  =>    DADOS_AUDIO <=  "0101111000111110";
						 when  28  =>    DADOS_AUDIO <=  "0110000011011010";
						 when  29  =>    DADOS_AUDIO <=  "0110001101011111";
						 when  30  =>    DADOS_AUDIO <=  "0110010111001100";
						 when  31  =>    DADOS_AUDIO <=  "0110100000100000";
						 when  32  =>    DADOS_AUDIO <=  "0110101001011100";
						 when  33  =>    DADOS_AUDIO <=  "0110110001111110";
						 when  34  =>    DADOS_AUDIO <=  "0110111010000101";
						 when  35  =>    DADOS_AUDIO <=  "0111000001110011";
						 when  36  =>    DADOS_AUDIO <=  "0111001001000101";
						 when  37  =>    DADOS_AUDIO <=  "0111001111111011";
						 when  38  =>    DADOS_AUDIO <=  "0111010110010110";
						 when  39  =>    DADOS_AUDIO <=  "0111011100010101";
						 when  40  =>    DADOS_AUDIO <=  "0111100001110111";
						 when  41  =>    DADOS_AUDIO <=  "0111100110111100";
						 when  42  =>    DADOS_AUDIO <=  "0111101011100011";
						 when  43  =>    DADOS_AUDIO <=  "0111101111101110";
						 when  44  =>    DADOS_AUDIO <=  "0111110011011010";
						 when  45  =>    DADOS_AUDIO <=  "0111110110101000";
						 when  46  =>    DADOS_AUDIO <=  "0111111001011000";
						 when  47  =>    DADOS_AUDIO <=  "0111111011101010";
						 when  48  =>    DADOS_AUDIO <=  "0111111101011101";
						 when  49  =>    DADOS_AUDIO <=  "0111111110110010";
						 when  50  =>    DADOS_AUDIO <=  "0111111111100111";
						 when  51  =>    DADOS_AUDIO <=  "0111111111111111";
						 when  52  =>    DADOS_AUDIO <=  "0111111111110111";
						 when  53  =>    DADOS_AUDIO <=  "0111111111010000";
						 when  54  =>    DADOS_AUDIO <=  "0111111110001011";
						 when  55  =>    DADOS_AUDIO <=  "0111111100100111";
						 when  56  =>    DADOS_AUDIO <=  "0111111010100101";
						 when  57  =>    DADOS_AUDIO <=  "0111111000000100";
						 when  58  =>    DADOS_AUDIO <=  "0111110101000101";
						 when  59  =>    DADOS_AUDIO <=  "0111110001100111";
						 when  60  =>    DADOS_AUDIO <=  "0111101101101100";
						 when  61  =>    DADOS_AUDIO <=  "0111101001010011";
						 when  62  =>    DADOS_AUDIO <=  "0111100100011101";
						 when  63  =>    DADOS_AUDIO <=  "0111011111001001";
						 when  64  =>    DADOS_AUDIO <=  "0111011001011001";
						 when  65  =>    DADOS_AUDIO <=  "0111010011001100";
						 when  66  =>    DADOS_AUDIO <=  "0111001100100100";
						 when  67  =>    DADOS_AUDIO <=  "0111000101011111";
						 when  68  =>    DADOS_AUDIO <=  "0110111101111111";
						 when  69  =>    DADOS_AUDIO <=  "0110110110000101";
						 when  70  =>    DADOS_AUDIO <=  "0110101101110000";
						 when  71  =>    DADOS_AUDIO <=  "0110100101000001";
						 when  72  =>    DADOS_AUDIO <=  "0110011011111001";
						 when  73  =>    DADOS_AUDIO <=  "0110010010011000";
						 when  74  =>    DADOS_AUDIO <=  "0110001000011111";
						 when  75  =>    DADOS_AUDIO <=  "0101111110001111";
						 when  76  =>    DADOS_AUDIO <=  "0101110011100111";
						 when  77  =>    DADOS_AUDIO <=  "0101101000101001";
						 when  78  =>    DADOS_AUDIO <=  "0101011101010101";
						 when  79  =>    DADOS_AUDIO <=  "0101010001101101";
						 when  80  =>    DADOS_AUDIO <=  "0101000101110000";
						 when  81  =>    DADOS_AUDIO <=  "0100111001011111";
						 when  82  =>    DADOS_AUDIO <=  "0100101100111100";
						 when  83  =>    DADOS_AUDIO <=  "0100100000000111";
						 when  84  =>    DADOS_AUDIO <=  "0100010011000000";
						 when  85  =>    DADOS_AUDIO <=  "0100000101101001";
						 when  86  =>    DADOS_AUDIO <=  "0011111000000010";
						 when  87  =>    DADOS_AUDIO <=  "0011101010001100";
						 when  88  =>    DADOS_AUDIO <=  "0011011100001000";
						 when  89  =>    DADOS_AUDIO <=  "0011001101110110";
						 when  90  =>    DADOS_AUDIO <=  "0010111111011001";
						 when  91  =>    DADOS_AUDIO <=  "0010110000110000";
						 when  92  =>    DADOS_AUDIO <=  "0010100001111100";
						 when  93  =>    DADOS_AUDIO <=  "0010010010111110";
						 when  94  =>    DADOS_AUDIO <=  "0010000011111000";
						 when  95  =>    DADOS_AUDIO <=  "0001110100101010";
						 when  96  =>    DADOS_AUDIO <=  "0001100101010101";
						 when  97  =>    DADOS_AUDIO <=  "0001010101111001";
						 when  98  =>    DADOS_AUDIO <=  "0001000110011001";
						 when  99  =>    DADOS_AUDIO <=  "0000110110110100";
						 when  100  =>    DADOS_AUDIO <=  "0000100111001100";
						 when  101  =>    DADOS_AUDIO <=  "0000010111100001";
						 when  102  =>    DADOS_AUDIO <=  "0000000111110110";
						 when  103  =>    DADOS_AUDIO <=  "1111111000001010";
						 when  104  =>    DADOS_AUDIO <=  "1111101000011111";
						 when  105  =>    DADOS_AUDIO <=  "1111011000110100";
						 when  106  =>    DADOS_AUDIO <=  "1111001001001100";
						 when  107  =>    DADOS_AUDIO <=  "1110111001100111";
						 when  108  =>    DADOS_AUDIO <=  "1110101010000111";
						 when  109  =>    DADOS_AUDIO <=  "1110011010101011";
						 when  110  =>    DADOS_AUDIO <=  "1110001011010110";
						 when  111  =>    DADOS_AUDIO <=  "1101111100001000";
						 when  112  =>    DADOS_AUDIO <=  "1101101101000010";
						 when  113  =>    DADOS_AUDIO <=  "1101011110000100";
						 when  114  =>    DADOS_AUDIO <=  "1101001111010000";
						 when  115  =>    DADOS_AUDIO <=  "1101000000100111";
						 when  116  =>    DADOS_AUDIO <=  "1100110010001010";
						 when  117  =>    DADOS_AUDIO <=  "1100100011111000";
						 when  118  =>    DADOS_AUDIO <=  "1100010101110100";
						 when  119  =>    DADOS_AUDIO <=  "1100000111111110";
						 when  120  =>    DADOS_AUDIO <=  "1011111010010111";
						 when  121  =>    DADOS_AUDIO <=  "1011101101000000";
						 when  122  =>    DADOS_AUDIO <=  "1011011111111001";
						 when  123  =>    DADOS_AUDIO <=  "1011010011000100";
						 when  124  =>    DADOS_AUDIO <=  "1011000110100001";
						 when  125  =>    DADOS_AUDIO <=  "1010111010010000";
						 when  126  =>    DADOS_AUDIO <=  "1010101110010011";
						 when  127  =>    DADOS_AUDIO <=  "1010100010101011";
						 when  128  =>    DADOS_AUDIO <=  "1010010111010111";
						 when  129  =>    DADOS_AUDIO <=  "1010001100011001";
						 when  130  =>    DADOS_AUDIO <=  "1010000001110001";
						 when  131  =>    DADOS_AUDIO <=  "1001110111100001";
						 when  132  =>    DADOS_AUDIO <=  "1001101101101000";
						 when  133  =>    DADOS_AUDIO <=  "1001100100000111";
						 when  134  =>    DADOS_AUDIO <=  "1001011010111111";
						 when  135  =>    DADOS_AUDIO <=  "1001010010010000";
						 when  136  =>    DADOS_AUDIO <=  "1001001001111011";
						 when  137  =>    DADOS_AUDIO <=  "1001000010000001";
						 when  138  =>    DADOS_AUDIO <=  "1000111010100001";
						 when  139  =>    DADOS_AUDIO <=  "1000110011011100";
						 when  140  =>    DADOS_AUDIO <=  "1000101100110100";
						 when  141  =>    DADOS_AUDIO <=  "1000100110100111";
						 when  142  =>    DADOS_AUDIO <=  "1000100000110111";
						 when  143  =>    DADOS_AUDIO <=  "1000011011100011";
						 when  144  =>    DADOS_AUDIO <=  "1000010110101101";
						 when  145  =>    DADOS_AUDIO <=  "1000010010010100";
						 when  146  =>    DADOS_AUDIO <=  "1000001110011001";
						 when  147  =>    DADOS_AUDIO <=  "1000001010111011";
						 when  148  =>    DADOS_AUDIO <=  "1000000111111100";
						 when  149  =>    DADOS_AUDIO <=  "1000000101011011";
						 when  150  =>    DADOS_AUDIO <=  "1000000011011001";
						 when  151  =>    DADOS_AUDIO <=  "1000000001110101";
						 when  152  =>    DADOS_AUDIO <=  "1000000000110000";
						 when  153  =>    DADOS_AUDIO <=  "1000000000001001";
						 when  154  =>    DADOS_AUDIO <=  "1000000000000001";
						 when  155  =>    DADOS_AUDIO <=  "1000000000011001";
						 when  156  =>    DADOS_AUDIO <=  "1000000001001110";
						 when  157  =>    DADOS_AUDIO <=  "1000000010100011";
						 when  158  =>    DADOS_AUDIO <=  "1000000100010110";
						 when  159  =>    DADOS_AUDIO <=  "1000000110101000";
						 when  160  =>    DADOS_AUDIO <=  "1000001001011000";
						 when  161  =>    DADOS_AUDIO <=  "1000001100100110";
						 when  162  =>    DADOS_AUDIO <=  "1000010000010010";
						 when  163  =>    DADOS_AUDIO <=  "1000010100011101";
						 when  164  =>    DADOS_AUDIO <=  "1000011001000100";
						 when  165  =>    DADOS_AUDIO <=  "1000011110001001";
						 when  166  =>    DADOS_AUDIO <=  "1000100011101011";
						 when  167  =>    DADOS_AUDIO <=  "1000101001101010";
						 when  168  =>    DADOS_AUDIO <=  "1000110000000101";
						 when  169  =>    DADOS_AUDIO <=  "1000110110111011";
						 when  170  =>    DADOS_AUDIO <=  "1000111110001101";
						 when  171  =>    DADOS_AUDIO <=  "1001000101111011";
						 when  172  =>    DADOS_AUDIO <=  "1001001110000010";
						 when  173  =>    DADOS_AUDIO <=  "1001010110100100";
						 when  174  =>    DADOS_AUDIO <=  "1001011111100000";
						 when  175  =>    DADOS_AUDIO <=  "1001101000110100";
						 when  176  =>    DADOS_AUDIO <=  "1001110010100001";
						 when  177  =>    DADOS_AUDIO <=  "1001111100100110";
						 when  178  =>    DADOS_AUDIO <=  "1010000111000010";
						 when  179  =>    DADOS_AUDIO <=  "1010010001110101";
						 when  180  =>    DADOS_AUDIO <=  "1010011100111110";
						 when  181  =>    DADOS_AUDIO <=  "1010101000011100";
						 when  182  =>    DADOS_AUDIO <=  "1010110100001111";
						 when  183  =>    DADOS_AUDIO <=  "1011000000010110";
						 when  184  =>    DADOS_AUDIO <=  "1011001100110000";
						 when  185  =>    DADOS_AUDIO <=  "1011011001011100";
						 when  186  =>    DADOS_AUDIO <=  "1011100110011011";
						 when  187  =>    DADOS_AUDIO <=  "1011110011101010";
						 when  188  =>    DADOS_AUDIO <=  "1100000001001001";
						 when  189  =>    DADOS_AUDIO <=  "1100001110111000";
						 when  190  =>    DADOS_AUDIO <=  "1100011100110101";
						 when  191  =>    DADOS_AUDIO <=  "1100101010111111";
						 when  192  =>    DADOS_AUDIO <=  "1100111001010111";
						 when  193  =>    DADOS_AUDIO <=  "1101000111111010";
						 when  194  =>    DADOS_AUDIO <=  "1101010110101001";
						 when  195  =>    DADOS_AUDIO <=  "1101100101100010";
						 when  196  =>    DADOS_AUDIO <=  "1101110100100100";
						 when  197  =>    DADOS_AUDIO <=  "1110000011101110";
						 when  198  =>    DADOS_AUDIO <=  "1110010011000000";
						 when  199  =>    DADOS_AUDIO <=  "1110100010011000";
						 when  200  =>    DADOS_AUDIO <=  "1110110001110110";
						 when  201  =>    DADOS_AUDIO <=  "1111000001011001";
						 when  202  =>    DADOS_AUDIO <=  "1111010001000000";
						 when  203  =>    DADOS_AUDIO <=  "1111100000101001";
						 when  204  =>    DADOS_AUDIO <=  "1111110000010100";
						 when  205  =>    DADOS_AUDIO <=  "0000000000000000";
						 when others =>	DADOS_AUDIO <=  "0000000000000000";
					end case;
				when 12 =>
					n_pontos <= 194;
					reset <= '0';
					case aux_dados is
					    when  0  =>    DADOS_AUDIO <=  "0000000000000000";
						 when  1  =>    DADOS_AUDIO <=  "0000010000101010";
						 when  2  =>    DADOS_AUDIO <=  "0000100001010100";
						 when  3  =>    DADOS_AUDIO <=  "0000110001111011";
						 when  4  =>    DADOS_AUDIO <=  "0001000010011111";
						 when  5  =>    DADOS_AUDIO <=  "0001010010111110";
						 when  6  =>    DADOS_AUDIO <=  "0001100011011000";
						 when  7  =>    DADOS_AUDIO <=  "0001110011101010";
						 when  8  =>    DADOS_AUDIO <=  "0010000011110110";
						 when  9  =>    DADOS_AUDIO <=  "0010010011111000";
						 when  10  =>    DADOS_AUDIO <=  "0010100011110000";
						 when  11  =>    DADOS_AUDIO <=  "0010110011011101";
						 when  12  =>    DADOS_AUDIO <=  "0011000010111110";
						 when  13  =>    DADOS_AUDIO <=  "0011010010010001";
						 when  14  =>    DADOS_AUDIO <=  "0011100001010111";
						 when  15  =>    DADOS_AUDIO <=  "0011110000001101";
						 when  16  =>    DADOS_AUDIO <=  "0011111110110010";
						 when  17  =>    DADOS_AUDIO <=  "0100001101000111";
						 when  18  =>    DADOS_AUDIO <=  "0100011011001001";
						 when  19  =>    DADOS_AUDIO <=  "0100101000111000";
						 when  20  =>    DADOS_AUDIO <=  "0100110110010011";
						 when  21  =>    DADOS_AUDIO <=  "0101000011011001";
						 when  22  =>    DADOS_AUDIO <=  "0101010000001001";
						 when  23  =>    DADOS_AUDIO <=  "0101011100100010";
						 when  24  =>    DADOS_AUDIO <=  "0101101000100011";
						 when  25  =>    DADOS_AUDIO <=  "0101110100001101";
						 when  26  =>    DADOS_AUDIO <=  "0101111111011100";
						 when  27  =>    DADOS_AUDIO <=  "0110001010010010";
						 when  28  =>    DADOS_AUDIO <=  "0110010100101101";
						 when  29  =>    DADOS_AUDIO <=  "0110011110101101";
						 when  30  =>    DADOS_AUDIO <=  "0110101000010000";
						 when  31  =>    DADOS_AUDIO <=  "0110110001010111";
						 when  32  =>    DADOS_AUDIO <=  "0110111010000000";
						 when  33  =>    DADOS_AUDIO <=  "0111000010001011";
						 when  34  =>    DADOS_AUDIO <=  "0111001001111000";
						 when  35  =>    DADOS_AUDIO <=  "0111010001000110";
						 when  36  =>    DADOS_AUDIO <=  "0111010111110100";
						 when  37  =>    DADOS_AUDIO <=  "0111011110000010";
						 when  38  =>    DADOS_AUDIO <=  "0111100011110000";
						 when  39  =>    DADOS_AUDIO <=  "0111101000111101";
						 when  40  =>    DADOS_AUDIO <=  "0111101101101001";
						 when  41  =>    DADOS_AUDIO <=  "0111110001110011";
						 when  42  =>    DADOS_AUDIO <=  "0111110101011100";
						 when  43  =>    DADOS_AUDIO <=  "0111111000100010";
						 when  44  =>    DADOS_AUDIO <=  "0111111011000110";
						 when  45  =>    DADOS_AUDIO <=  "0111111101001000";
						 when  46  =>    DADOS_AUDIO <=  "0111111110101000";
						 when  47  =>    DADOS_AUDIO <=  "0111111111100100";
						 when  48  =>    DADOS_AUDIO <=  "0111111111111110";
						 when  49  =>    DADOS_AUDIO <=  "0111111111110110";
						 when  50  =>    DADOS_AUDIO <=  "0111111111001010";
						 when  51  =>    DADOS_AUDIO <=  "0111111101111100";
						 when  52  =>    DADOS_AUDIO <=  "0111111100001100";
						 when  53  =>    DADOS_AUDIO <=  "0111111001111000";
						 when  54  =>    DADOS_AUDIO <=  "0111110111000011";
						 when  55  =>    DADOS_AUDIO <=  "0111110011101100";
						 when  56  =>    DADOS_AUDIO <=  "0111101111110010";
						 when  57  =>    DADOS_AUDIO <=  "0111101011010111";
						 when  58  =>    DADOS_AUDIO <=  "0111100110011011";
						 when  59  =>    DADOS_AUDIO <=  "0111100000111101";
						 when  60  =>    DADOS_AUDIO <=  "0111011010111111";
						 when  61  =>    DADOS_AUDIO <=  "0111010100100001";
						 when  62  =>    DADOS_AUDIO <=  "0111001101100011";
						 when  63  =>    DADOS_AUDIO <=  "0111000110000110";
						 when  64  =>    DADOS_AUDIO <=  "0110111110001010";
						 when  65  =>    DADOS_AUDIO <=  "0110110101101111";
						 when  66  =>    DADOS_AUDIO <=  "0110101100110111";
						 when  67  =>    DADOS_AUDIO <=  "0110100011100010";
						 when  68  =>    DADOS_AUDIO <=  "0110011001110000";
						 when  69  =>    DADOS_AUDIO <=  "0110001111100011";
						 when  70  =>    DADOS_AUDIO <=  "0110000100111010";
						 when  71  =>    DADOS_AUDIO <=  "0101111001111000";
						 when  72  =>    DADOS_AUDIO <=  "0101101110011011";
						 when  73  =>    DADOS_AUDIO <=  "0101100010100110";
						 when  74  =>    DADOS_AUDIO <=  "0101010110011000";
						 when  75  =>    DADOS_AUDIO <=  "0101001001110100";
						 when  76  =>    DADOS_AUDIO <=  "0100111100111001";
						 when  77  =>    DADOS_AUDIO <=  "0100101111101000";
						 when  78  =>    DADOS_AUDIO <=  "0100100010000011";
						 when  79  =>    DADOS_AUDIO <=  "0100010100001010";
						 when  80  =>    DADOS_AUDIO <=  "0100000101111111";
						 when  81  =>    DADOS_AUDIO <=  "0011110111100010";
						 when  82  =>    DADOS_AUDIO <=  "0011101000110100";
						 when  83  =>    DADOS_AUDIO <=  "0011011001110110";
						 when  84  =>    DADOS_AUDIO <=  "0011001010101001";
						 when  85  =>    DADOS_AUDIO <=  "0010111011001111";
						 when  86  =>    DADOS_AUDIO <=  "0010101011101000";
						 when  87  =>    DADOS_AUDIO <=  "0010011011110101";
						 when  88  =>    DADOS_AUDIO <=  "0010001011111000";
						 when  89  =>    DADOS_AUDIO <=  "0001111011110001";
						 when  90  =>    DADOS_AUDIO <=  "0001101011100010";
						 when  91  =>    DADOS_AUDIO <=  "0001011011001011";
						 when  92  =>    DADOS_AUDIO <=  "0001001010101111";
						 when  93  =>    DADOS_AUDIO <=  "0000111010001101";
						 when  94  =>    DADOS_AUDIO <=  "0000101001100111";
						 when  95  =>    DADOS_AUDIO <=  "0000011000111111";
						 when  96  =>    DADOS_AUDIO <=  "0000001000010101";
						 when  97  =>    DADOS_AUDIO <=  "1111110111101011";
						 when  98  =>    DADOS_AUDIO <=  "1111100111000001";
						 when  99  =>    DADOS_AUDIO <=  "1111010110011001";
						 when  100  =>    DADOS_AUDIO <=  "1111000101110011";
						 when  101  =>    DADOS_AUDIO <=  "1110110101010001";
						 when  102  =>    DADOS_AUDIO <=  "1110100100110101";
						 when  103  =>    DADOS_AUDIO <=  "1110010100011110";
						 when  104  =>    DADOS_AUDIO <=  "1110000100001111";
						 when  105  =>    DADOS_AUDIO <=  "1101110100001000";
						 when  106  =>    DADOS_AUDIO <=  "1101100100001011";
						 when  107  =>    DADOS_AUDIO <=  "1101010100011000";
						 when  108  =>    DADOS_AUDIO <=  "1101000100110001";
						 when  109  =>    DADOS_AUDIO <=  "1100110101010111";
						 when  110  =>    DADOS_AUDIO <=  "1100100110001010";
						 when  111  =>    DADOS_AUDIO <=  "1100010111001100";
						 when  112  =>    DADOS_AUDIO <=  "1100001000011110";
						 when  113  =>    DADOS_AUDIO <=  "1011111010000001";
						 when  114  =>    DADOS_AUDIO <=  "1011101011110110";
						 when  115  =>    DADOS_AUDIO <=  "1011011101111101";
						 when  116  =>    DADOS_AUDIO <=  "1011010000011000";
						 when  117  =>    DADOS_AUDIO <=  "1011000011000111";
						 when  118  =>    DADOS_AUDIO <=  "1010110110001100";
						 when  119  =>    DADOS_AUDIO <=  "1010101001101000";
						 when  120  =>    DADOS_AUDIO <=  "1010011101011010";
						 when  121  =>    DADOS_AUDIO <=  "1010010001100101";
						 when  122  =>    DADOS_AUDIO <=  "1010000110001000";
						 when  123  =>    DADOS_AUDIO <=  "1001111011000110";
						 when  124  =>    DADOS_AUDIO <=  "1001110000011101";
						 when  125  =>    DADOS_AUDIO <=  "1001100110010000";
						 when  126  =>    DADOS_AUDIO <=  "1001011100011110";
						 when  127  =>    DADOS_AUDIO <=  "1001010011001001";
						 when  128  =>    DADOS_AUDIO <=  "1001001010010001";
						 when  129  =>    DADOS_AUDIO <=  "1001000001110110";
						 when  130  =>    DADOS_AUDIO <=  "1000111001111010";
						 when  131  =>    DADOS_AUDIO <=  "1000110010011101";
						 when  132  =>    DADOS_AUDIO <=  "1000101011011111";
						 when  133  =>    DADOS_AUDIO <=  "1000100101000001";
						 when  134  =>    DADOS_AUDIO <=  "1000011111000011";
						 when  135  =>    DADOS_AUDIO <=  "1000011001100101";
						 when  136  =>    DADOS_AUDIO <=  "1000010100101001";
						 when  137  =>    DADOS_AUDIO <=  "1000010000001110";
						 when  138  =>    DADOS_AUDIO <=  "1000001100010100";
						 when  139  =>    DADOS_AUDIO <=  "1000001000111101";
						 when  140  =>    DADOS_AUDIO <=  "1000000110001000";
						 when  141  =>    DADOS_AUDIO <=  "1000000011110100";
						 when  142  =>    DADOS_AUDIO <=  "1000000010000100";
						 when  143  =>    DADOS_AUDIO <=  "1000000000110110";
						 when  144  =>    DADOS_AUDIO <=  "1000000000001010";
						 when  145  =>    DADOS_AUDIO <=  "1000000000000010";
						 when  146  =>    DADOS_AUDIO <=  "1000000000011100";
						 when  147  =>    DADOS_AUDIO <=  "1000000001011000";
						 when  148  =>    DADOS_AUDIO <=  "1000000010111000";
						 when  149  =>    DADOS_AUDIO <=  "1000000100111010";
						 when  150  =>    DADOS_AUDIO <=  "1000000111011110";
						 when  151  =>    DADOS_AUDIO <=  "1000001010100100";
						 when  152  =>    DADOS_AUDIO <=  "1000001110001101";
						 when  153  =>    DADOS_AUDIO <=  "1000010010010111";
						 when  154  =>    DADOS_AUDIO <=  "1000010111000011";
						 when  155  =>    DADOS_AUDIO <=  "1000011100010000";
						 when  156  =>    DADOS_AUDIO <=  "1000100001111110";
						 when  157  =>    DADOS_AUDIO <=  "1000101000001100";
						 when  158  =>    DADOS_AUDIO <=  "1000101110111010";
						 when  159  =>    DADOS_AUDIO <=  "1000110110001000";
						 when  160  =>    DADOS_AUDIO <=  "1000111101110101";
						 when  161  =>    DADOS_AUDIO <=  "1001000110000000";
						 when  162  =>    DADOS_AUDIO <=  "1001001110101001";
						 when  163  =>    DADOS_AUDIO <=  "1001010111110000";
						 when  164  =>    DADOS_AUDIO <=  "1001100001010011";
						 when  165  =>    DADOS_AUDIO <=  "1001101011010011";
						 when  166  =>    DADOS_AUDIO <=  "1001110101101110";
						 when  167  =>    DADOS_AUDIO <=  "1010000000100100";
						 when  168  =>    DADOS_AUDIO <=  "1010001011110011";
						 when  169  =>    DADOS_AUDIO <=  "1010010111011101";
						 when  170  =>    DADOS_AUDIO <=  "1010100011011110";
						 when  171  =>    DADOS_AUDIO <=  "1010101111110111";
						 when  172  =>    DADOS_AUDIO <=  "1010111100100111";
						 when  173  =>    DADOS_AUDIO <=  "1011001001101101";
						 when  174  =>    DADOS_AUDIO <=  "1011010111001000";
						 when  175  =>    DADOS_AUDIO <=  "1011100100110111";
						 when  176  =>    DADOS_AUDIO <=  "1011110010111001";
						 when  177  =>    DADOS_AUDIO <=  "1100000001001110";
						 when  178  =>    DADOS_AUDIO <=  "1100001111110011";
						 when  179  =>    DADOS_AUDIO <=  "1100011110101001";
						 when  180  =>    DADOS_AUDIO <=  "1100101101101111";
						 when  181  =>    DADOS_AUDIO <=  "1100111101000010";
						 when  182  =>    DADOS_AUDIO <=  "1101001100100011";
						 when  183  =>    DADOS_AUDIO <=  "1101011100010000";
						 when  184  =>    DADOS_AUDIO <=  "1101101100001000";
						 when  185  =>    DADOS_AUDIO <=  "1101111100001010";
						 when  186  =>    DADOS_AUDIO <=  "1110001100010110";
						 when  187  =>    DADOS_AUDIO <=  "1110011100101000";
						 when  188  =>    DADOS_AUDIO <=  "1110101101000010";
						 when  189  =>    DADOS_AUDIO <=  "1110111101100001";
						 when  190  =>    DADOS_AUDIO <=  "1111001110000101";
						 when  191  =>    DADOS_AUDIO <=  "1111011110101100";
						 when  192  =>    DADOS_AUDIO <=  "1111101111010110";
						 when  193  =>    DADOS_AUDIO <=  "0000000000000000";
						 when others =>	DADOS_AUDIO <=  "0000000000000000";
					end case;
				when others =>
					reset <= '1';
			end case;
		end process;
	
			
end behavior;